// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire net76;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net77;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net78;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net114;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net115;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net116;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net144;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net145;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net146;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net147;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net148;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net149;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire \mod.buffer[0] ;
 wire \mod.buffer[100] ;
 wire \mod.buffer[101] ;
 wire \mod.buffer[102] ;
 wire \mod.buffer[103] ;
 wire \mod.buffer[104] ;
 wire \mod.buffer[105] ;
 wire \mod.buffer[106] ;
 wire \mod.buffer[107] ;
 wire \mod.buffer[108] ;
 wire \mod.buffer[109] ;
 wire \mod.buffer[10] ;
 wire \mod.buffer[110] ;
 wire \mod.buffer[111] ;
 wire \mod.buffer[112] ;
 wire \mod.buffer[113] ;
 wire \mod.buffer[114] ;
 wire \mod.buffer[115] ;
 wire \mod.buffer[116] ;
 wire \mod.buffer[117] ;
 wire \mod.buffer[118] ;
 wire \mod.buffer[119] ;
 wire \mod.buffer[11] ;
 wire \mod.buffer[120] ;
 wire \mod.buffer[121] ;
 wire \mod.buffer[122] ;
 wire \mod.buffer[123] ;
 wire \mod.buffer[124] ;
 wire \mod.buffer[125] ;
 wire \mod.buffer[126] ;
 wire \mod.buffer[127] ;
 wire \mod.buffer[128] ;
 wire \mod.buffer[129] ;
 wire \mod.buffer[12] ;
 wire \mod.buffer[130] ;
 wire \mod.buffer[131] ;
 wire \mod.buffer[132] ;
 wire \mod.buffer[133] ;
 wire \mod.buffer[134] ;
 wire \mod.buffer[135] ;
 wire \mod.buffer[136] ;
 wire \mod.buffer[137] ;
 wire \mod.buffer[138] ;
 wire \mod.buffer[139] ;
 wire \mod.buffer[13] ;
 wire \mod.buffer[14] ;
 wire \mod.buffer[15] ;
 wire \mod.buffer[16] ;
 wire \mod.buffer[17] ;
 wire \mod.buffer[18] ;
 wire \mod.buffer[19] ;
 wire \mod.buffer[1] ;
 wire \mod.buffer[20] ;
 wire \mod.buffer[21] ;
 wire \mod.buffer[22] ;
 wire \mod.buffer[23] ;
 wire \mod.buffer[24] ;
 wire \mod.buffer[25] ;
 wire \mod.buffer[26] ;
 wire \mod.buffer[27] ;
 wire \mod.buffer[28] ;
 wire \mod.buffer[29] ;
 wire \mod.buffer[2] ;
 wire \mod.buffer[30] ;
 wire \mod.buffer[31] ;
 wire \mod.buffer[32] ;
 wire \mod.buffer[33] ;
 wire \mod.buffer[34] ;
 wire \mod.buffer[35] ;
 wire \mod.buffer[36] ;
 wire \mod.buffer[37] ;
 wire \mod.buffer[38] ;
 wire \mod.buffer[39] ;
 wire \mod.buffer[3] ;
 wire \mod.buffer[40] ;
 wire \mod.buffer[41] ;
 wire \mod.buffer[42] ;
 wire \mod.buffer[43] ;
 wire \mod.buffer[44] ;
 wire \mod.buffer[45] ;
 wire \mod.buffer[46] ;
 wire \mod.buffer[47] ;
 wire \mod.buffer[48] ;
 wire \mod.buffer[49] ;
 wire \mod.buffer[4] ;
 wire \mod.buffer[50] ;
 wire \mod.buffer[51] ;
 wire \mod.buffer[52] ;
 wire \mod.buffer[53] ;
 wire \mod.buffer[54] ;
 wire \mod.buffer[55] ;
 wire \mod.buffer[56] ;
 wire \mod.buffer[57] ;
 wire \mod.buffer[58] ;
 wire \mod.buffer[59] ;
 wire \mod.buffer[5] ;
 wire \mod.buffer[60] ;
 wire \mod.buffer[61] ;
 wire \mod.buffer[62] ;
 wire \mod.buffer[63] ;
 wire \mod.buffer[64] ;
 wire \mod.buffer[65] ;
 wire \mod.buffer[66] ;
 wire \mod.buffer[67] ;
 wire \mod.buffer[68] ;
 wire \mod.buffer[69] ;
 wire \mod.buffer[6] ;
 wire \mod.buffer[70] ;
 wire \mod.buffer[71] ;
 wire \mod.buffer[72] ;
 wire \mod.buffer[73] ;
 wire \mod.buffer[74] ;
 wire \mod.buffer[75] ;
 wire \mod.buffer[76] ;
 wire \mod.buffer[77] ;
 wire \mod.buffer[78] ;
 wire \mod.buffer[79] ;
 wire \mod.buffer[7] ;
 wire \mod.buffer[80] ;
 wire \mod.buffer[81] ;
 wire \mod.buffer[82] ;
 wire \mod.buffer[83] ;
 wire \mod.buffer[84] ;
 wire \mod.buffer[85] ;
 wire \mod.buffer[86] ;
 wire \mod.buffer[87] ;
 wire \mod.buffer[88] ;
 wire \mod.buffer[89] ;
 wire \mod.buffer[8] ;
 wire \mod.buffer[90] ;
 wire \mod.buffer[91] ;
 wire \mod.buffer[92] ;
 wire \mod.buffer[93] ;
 wire \mod.buffer[94] ;
 wire \mod.buffer[95] ;
 wire \mod.buffer[96] ;
 wire \mod.buffer[97] ;
 wire \mod.buffer[98] ;
 wire \mod.buffer[99] ;
 wire \mod.buffer[9] ;
 wire \mod.counter[0] ;
 wire \mod.counter[1] ;
 wire \mod.counter[2] ;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net213;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net214;
 wire net242;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0881_ (.I(\mod.counter[0] ),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0882_ (.I(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0883_ (.I(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0884_ (.I(_0254_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0885_ (.A1(net1),
    .A2(\mod.buffer[6] ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0886_ (.A1(_0255_),
    .A2(_0256_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0887_ (.I(\mod.counter[1] ),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0888_ (.A1(_0257_),
    .A2(\mod.counter[0] ),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0889_ (.I(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0890_ (.A1(_0256_),
    .A2(_0259_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0891_ (.I(_0252_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0892_ (.I(\mod.counter[2] ),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0893_ (.I(_0261_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0894_ (.A1(_0260_),
    .A2(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0895_ (.I(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0896_ (.I(\mod.counter[1] ),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0897_ (.I(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0898_ (.I(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0899_ (.A1(_0266_),
    .A2(_0253_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0900_ (.I(\mod.counter[2] ),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0901_ (.I(_0269_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0902_ (.I0(_0267_),
    .I1(_0268_),
    .S(_0270_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0903_ (.A1(_0264_),
    .A2(_0271_),
    .B(_0256_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0904_ (.I(\mod.buffer[6] ),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0905_ (.I(\mod.buffer[5] ),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0906_ (.A1(_0272_),
    .A2(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0907_ (.I(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0908_ (.I(\mod.buffer[1] ),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0909_ (.I(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0910_ (.I(_0277_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0911_ (.I(\mod.buffer[0] ),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0912_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0913_ (.I(_0265_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0914_ (.I(\mod.counter[2] ),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0915_ (.A1(_0281_),
    .A2(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0916_ (.I(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0917_ (.I(\mod.counter[0] ),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0918_ (.A1(_0281_),
    .A2(_0285_),
    .A3(_0282_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0919_ (.I(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0920_ (.A1(_0280_),
    .A2(_0284_),
    .A3(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0921_ (.I(\mod.buffer[0] ),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0922_ (.I(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0923_ (.I(\mod.buffer[1] ),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0924_ (.I(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0925_ (.A1(_0290_),
    .A2(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0926_ (.I(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0927_ (.A1(_0267_),
    .A2(_0254_),
    .A3(_0270_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0928_ (.I(_0265_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0929_ (.I(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0930_ (.I(_0262_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0931_ (.A1(_0297_),
    .A2(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0932_ (.A1(_0295_),
    .A2(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0933_ (.I(\mod.buffer[2] ),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0934_ (.I(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _0935_ (.A1(_0278_),
    .A2(_0288_),
    .B1(_0294_),
    .B2(_0300_),
    .C(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0936_ (.I(_0289_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0937_ (.I(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0938_ (.A1(_0265_),
    .A2(_0261_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0939_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0940_ (.I(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0941_ (.A1(_0305_),
    .A2(_0259_),
    .B(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0942_ (.I(_0276_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0943_ (.A1(_0310_),
    .A2(_0301_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0944_ (.I(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0945_ (.I(\mod.buffer[2] ),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0946_ (.A1(_0257_),
    .A2(_0252_),
    .A3(\mod.counter[2] ),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0947_ (.A1(_0290_),
    .A2(_0314_),
    .A3(_0286_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0948_ (.I(_0282_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0949_ (.A1(_0266_),
    .A2(_0285_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0950_ (.A1(_0316_),
    .A2(_0317_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0951_ (.A1(_0316_),
    .A2(_0317_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0952_ (.I(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0953_ (.A1(_0313_),
    .A2(_0315_),
    .A3(_0318_),
    .A4(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0954_ (.I(_0285_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0955_ (.A1(_0322_),
    .A2(_0284_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0956_ (.I(\mod.buffer[0] ),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0957_ (.I(_0324_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0958_ (.A1(_0325_),
    .A2(_0287_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0959_ (.A1(_0323_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0960_ (.A1(_0305_),
    .A2(_0271_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0961_ (.I(_0310_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0962_ (.I(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0963_ (.A1(_0312_),
    .A2(_0321_),
    .B1(_0328_),
    .B2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0964_ (.I(\mod.buffer[3] ),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0965_ (.I(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0966_ (.A1(_0303_),
    .A2(_0309_),
    .B(_0331_),
    .C(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0967_ (.I(\mod.buffer[4] ),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0968_ (.I(_0301_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0969_ (.I(_0257_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0970_ (.I(_0269_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0971_ (.A1(_0337_),
    .A2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0972_ (.A1(_0339_),
    .A2(_0319_),
    .B(_0304_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0973_ (.I(_0296_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0974_ (.I(_0252_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0975_ (.A1(_0341_),
    .A2(_0342_),
    .A3(_0338_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0976_ (.I(_0260_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0977_ (.A1(_0344_),
    .A2(_0283_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0978_ (.I(_0324_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0979_ (.A1(_0343_),
    .A2(_0345_),
    .B(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0980_ (.I(_0276_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0981_ (.I(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0982_ (.I(\mod.buffer[2] ),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0983_ (.I(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0984_ (.A1(_0349_),
    .A2(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0985_ (.A1(_0336_),
    .A2(_0340_),
    .A3(_0347_),
    .B(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0986_ (.A1(_0341_),
    .A2(_0322_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0987_ (.A1(_0281_),
    .A2(_0260_),
    .A3(_0282_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0988_ (.I(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0989_ (.A1(_0354_),
    .A2(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0990_ (.I(_0289_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0991_ (.A1(_0358_),
    .A2(_0310_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0992_ (.A1(_0263_),
    .A2(_0299_),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0993_ (.A1(_0294_),
    .A2(_0357_),
    .B(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0994_ (.I(_0276_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0995_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0996_ (.I(_0260_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0997_ (.A1(_0364_),
    .A2(_0298_),
    .B(_0267_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0998_ (.I(_0290_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0999_ (.A1(_0343_),
    .A2(_0365_),
    .B(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1000_ (.A1(_0280_),
    .A2(_0318_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1001_ (.I(_0348_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1002_ (.I(_0306_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1003_ (.A1(_0346_),
    .A2(_0258_),
    .A3(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1004_ (.A1(_0369_),
    .A2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1005_ (.A1(_0337_),
    .A2(_0344_),
    .A3(_0298_),
    .A4(_0325_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1006_ (.A1(_0296_),
    .A2(_0342_),
    .A3(_0324_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1007_ (.I(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _1008_ (.A1(_0363_),
    .A2(_0367_),
    .A3(_0368_),
    .B1(_0372_),
    .B2(_0373_),
    .B3(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1009_ (.I(\mod.buffer[2] ),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1010_ (.I(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1011_ (.I(\mod.buffer[3] ),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1012_ (.I(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1013_ (.A1(_0353_),
    .A2(_0361_),
    .B1(_0376_),
    .B2(_0378_),
    .C(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1014_ (.A1(_0335_),
    .A2(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1015_ (.I(\mod.buffer[0] ),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1016_ (.A1(_0253_),
    .A2(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1017_ (.A1(_0341_),
    .A2(_0269_),
    .A3(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1018_ (.I(_0261_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1019_ (.A1(_0266_),
    .A2(_0344_),
    .A3(_0386_),
    .A4(_0279_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1020_ (.A1(_0385_),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1021_ (.I(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1022_ (.I(_0291_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1023_ (.I(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1024_ (.A1(_0326_),
    .A2(_0389_),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1025_ (.I(_0350_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1026_ (.A1(_0364_),
    .A2(_0390_),
    .A3(_0370_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1027_ (.A1(_0393_),
    .A2(_0394_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1028_ (.I(_0383_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1029_ (.I(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1030_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1031_ (.I(_0313_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1032_ (.A1(_0398_),
    .A2(_0308_),
    .B(_0288_),
    .C(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1033_ (.I(\mod.buffer[3] ),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1034_ (.I(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1035_ (.A1(_0392_),
    .A2(_0395_),
    .B(_0400_),
    .C(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1036_ (.I(\mod.buffer[4] ),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1037_ (.I(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1038_ (.I(_0363_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1039_ (.I(_0343_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1040_ (.A1(_0323_),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1041_ (.A1(_0313_),
    .A2(_0379_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1042_ (.I(_0310_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1043_ (.A1(_0397_),
    .A2(_0287_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1044_ (.A1(_0406_),
    .A2(_0408_),
    .B(_0409_),
    .C(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1045_ (.A1(_0405_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1046_ (.A1(_0334_),
    .A2(_0382_),
    .B1(_0403_),
    .B2(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1047_ (.I(_0272_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1048_ (.A1(_0415_),
    .A2(net4),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1049_ (.I(\mod.buffer[3] ),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1050_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1051_ (.I(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1052_ (.I(_0352_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1053_ (.I(_0359_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1054_ (.A1(_0348_),
    .A2(_0350_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1055_ (.I(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1056_ (.I(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1057_ (.A1(_0308_),
    .A2(_0420_),
    .A3(_0421_),
    .A4(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1058_ (.I(_0351_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1059_ (.A1(_0426_),
    .A2(_0401_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1060_ (.A1(_0386_),
    .A2(_0268_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1061_ (.I(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1062_ (.A1(_0257_),
    .A2(_0261_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1063_ (.A1(_0279_),
    .A2(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1064_ (.I(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1065_ (.I(_0292_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1066_ (.A1(_0433_),
    .A2(_0430_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1067_ (.A1(_0401_),
    .A2(_0429_),
    .A3(_0432_),
    .A4(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1068_ (.A1(_0427_),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1069_ (.I(_0315_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1070_ (.A1(_0290_),
    .A2(_0306_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1071_ (.I(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1072_ (.A1(_0329_),
    .A2(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1073_ (.I(_0322_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1074_ (.I(_0351_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1075_ (.A1(_0271_),
    .A2(_0437_),
    .B1(_0440_),
    .B2(_0441_),
    .C(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1076_ (.A1(_0436_),
    .A2(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1077_ (.I(\mod.buffer[4] ),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1078_ (.I(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1079_ (.A1(_0419_),
    .A2(_0425_),
    .B(_0444_),
    .C(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1080_ (.A1(_0281_),
    .A2(_0285_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1081_ (.I(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1082_ (.A1(_0449_),
    .A2(_0434_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1083_ (.A1(_0358_),
    .A2(_0362_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1084_ (.A1(_0428_),
    .A2(_0451_),
    .B(_0377_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1085_ (.A1(_0429_),
    .A2(_0294_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1086_ (.I(_0302_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1087_ (.I(_0445_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1088_ (.A1(_0380_),
    .A2(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1089_ (.A1(_0450_),
    .A2(_0452_),
    .B1(_0453_),
    .B2(_0454_),
    .C(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1090_ (.A1(_0415_),
    .A2(_0273_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1091_ (.A1(_0447_),
    .A2(_0457_),
    .B(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1092_ (.A1(_0275_),
    .A2(_0414_),
    .B(_0416_),
    .C(_0459_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1093_ (.I(_0272_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1094_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1095_ (.I(_0305_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1096_ (.I(_0301_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1097_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1098_ (.I(_0390_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1099_ (.A1(_0396_),
    .A2(_0306_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1100_ (.A1(_0259_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1101_ (.A1(_0254_),
    .A2(_0270_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1102_ (.I(_0345_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1103_ (.I(_0279_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1104_ (.A1(_0468_),
    .A2(_0469_),
    .B(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1105_ (.I(_0384_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1106_ (.I(_0348_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1107_ (.A1(_0297_),
    .A2(_0322_),
    .A3(_0316_),
    .A4(_0396_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1108_ (.A1(_0473_),
    .A2(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1109_ (.A1(_0465_),
    .A2(_0467_),
    .A3(_0471_),
    .B1(_0472_),
    .B2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1110_ (.A1(_0464_),
    .A2(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1111_ (.I(_0410_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1112_ (.I(_0338_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1113_ (.I(_0346_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1114_ (.A1(_0341_),
    .A2(_0342_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1115_ (.I(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1116_ (.A1(_0397_),
    .A2(_0449_),
    .A3(_0307_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1117_ (.A1(_0479_),
    .A2(_0480_),
    .A3(_0482_),
    .B(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1118_ (.A1(_0344_),
    .A2(_0283_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1119_ (.A1(_0355_),
    .A2(_0485_),
    .B(_0358_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1120_ (.A1(_0325_),
    .A2(_0428_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1121_ (.I(_0487_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1122_ (.I(_0277_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1123_ (.A1(_0486_),
    .A2(_0488_),
    .B(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1124_ (.A1(_0478_),
    .A2(_0484_),
    .B(_0490_),
    .C(_0464_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1125_ (.I(_0332_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1126_ (.A1(_0477_),
    .A2(_0491_),
    .B(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1127_ (.I(_0354_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1128_ (.I(_0486_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1129_ (.A1(_0442_),
    .A2(_0495_),
    .A3(_0483_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1130_ (.A1(_0448_),
    .A2(_0431_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1131_ (.A1(_0470_),
    .A2(_0354_),
    .B(_0351_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1132_ (.I(_0277_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1133_ (.A1(_0497_),
    .A2(_0498_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1134_ (.I(_0417_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1135_ (.A1(_0478_),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0500_),
    .C(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1136_ (.A1(_0405_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1137_ (.A1(_0433_),
    .A2(_0347_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1138_ (.A1(_0478_),
    .A2(_0494_),
    .B(_0409_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1139_ (.A1(_0479_),
    .A2(_0448_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1140_ (.A1(_0262_),
    .A2(_0383_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1141_ (.A1(_0296_),
    .A2(_0342_),
    .A3(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1142_ (.I(_0508_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1143_ (.A1(_0366_),
    .A2(_0506_),
    .B(_0509_),
    .C(_0356_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1144_ (.A1(_0499_),
    .A2(_0510_),
    .B(_0395_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1145_ (.A1(_0378_),
    .A2(_0375_),
    .A3(_0389_),
    .B(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1146_ (.A1(_0504_),
    .A2(_0505_),
    .B1(_0512_),
    .B2(_0492_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1147_ (.I(\mod.buffer[4] ),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1148_ (.A1(_0493_),
    .A2(_0503_),
    .B1(_0513_),
    .B2(_0514_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1149_ (.I(\mod.buffer[5] ),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1150_ (.A1(_0272_),
    .A2(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1151_ (.I(_0473_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1152_ (.A1(_0253_),
    .A2(_0383_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1153_ (.A1(_0337_),
    .A2(_0386_),
    .A3(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1154_ (.I(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1155_ (.A1(_0521_),
    .A2(_0509_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1156_ (.A1(_0270_),
    .A2(_0304_),
    .A3(_0354_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1157_ (.A1(_0518_),
    .A2(_0399_),
    .A3(_0522_),
    .A4(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1158_ (.I(_0485_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1159_ (.A1(_0356_),
    .A2(_0525_),
    .B(_0410_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1160_ (.A1(_0337_),
    .A2(_0338_),
    .A3(_0396_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1161_ (.A1(_0349_),
    .A2(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1162_ (.A1(_0463_),
    .A2(_0347_),
    .A3(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1163_ (.A1(_0259_),
    .A2(_0431_),
    .B(_0521_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1164_ (.I(_0422_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1165_ (.A1(_0526_),
    .A2(_0529_),
    .B1(_0530_),
    .B2(_0531_),
    .C(_0332_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1166_ (.I(_0311_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1167_ (.A1(_0433_),
    .A2(_0393_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1168_ (.I(_0356_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1169_ (.A1(_0535_),
    .A2(_0525_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1170_ (.A1(_0390_),
    .A2(_0313_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1171_ (.A1(_0428_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1172_ (.A1(_0533_),
    .A2(_0522_),
    .B1(_0534_),
    .B2(_0536_),
    .C(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1173_ (.I(_0417_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1174_ (.A1(_0524_),
    .A2(_0532_),
    .B1(_0539_),
    .B2(_0540_),
    .C(_0455_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1175_ (.A1(_0357_),
    .A2(_0451_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1176_ (.A1(_0464_),
    .A2(_0453_),
    .A3(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1177_ (.I(_0393_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1178_ (.A1(_0465_),
    .A2(_0340_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1179_ (.A1(_0544_),
    .A2(_0450_),
    .A3(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1180_ (.A1(_0543_),
    .A2(_0546_),
    .B(_0456_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1181_ (.A1(_0346_),
    .A2(_0362_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1182_ (.A1(_0548_),
    .A2(_0469_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1183_ (.A1(_0418_),
    .A2(_0455_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1184_ (.I(_0487_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1185_ (.A1(_0352_),
    .A2(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1186_ (.A1(_0454_),
    .A2(_0549_),
    .B(_0550_),
    .C(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1187_ (.A1(_0517_),
    .A2(_0541_),
    .A3(_0547_),
    .A4(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1188_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0275_),
    .B2(_0515_),
    .C(_0554_),
    .ZN(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1189_ (.I(_0465_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1190_ (.A1(_0482_),
    .A2(_0469_),
    .B(_0397_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1191_ (.I(_0316_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1192_ (.A1(_0557_),
    .A2(_0519_),
    .B(_0391_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1193_ (.A1(_0391_),
    .A2(_0525_),
    .B1(_0556_),
    .B2(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1194_ (.I(_0349_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1195_ (.A1(_0297_),
    .A2(_0557_),
    .A3(_0472_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1196_ (.A1(_0560_),
    .A2(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1197_ (.A1(_0358_),
    .A2(_0284_),
    .A3(_0287_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1198_ (.A1(_0369_),
    .A2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1199_ (.A1(_0441_),
    .A2(_0439_),
    .B(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1200_ (.I(_0377_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1201_ (.A1(_0373_),
    .A2(_0562_),
    .B(_0565_),
    .C(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1202_ (.I(_0379_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1203_ (.A1(_0454_),
    .A2(_0559_),
    .B(_0567_),
    .C(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1204_ (.I(_0463_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1205_ (.A1(_0536_),
    .A2(_0534_),
    .B(_0538_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1206_ (.A1(_0570_),
    .A2(_0549_),
    .B(_0571_),
    .C(_0380_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1207_ (.A1(_0446_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1208_ (.A1(_0420_),
    .A2(_0551_),
    .B1(_0561_),
    .B2(_0312_),
    .C(_0402_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1209_ (.A1(_0437_),
    .A2(_0497_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1210_ (.A1(_0537_),
    .A2(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1211_ (.A1(_0369_),
    .A2(_0377_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1212_ (.A1(_0441_),
    .A2(_0426_),
    .A3(_0339_),
    .B1(_0423_),
    .B2(_0482_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1213_ (.A1(_0340_),
    .A2(_0577_),
    .B1(_0578_),
    .B2(_0398_),
    .C(_0501_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1214_ (.A1(_0576_),
    .A2(_0579_),
    .B(_0335_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1215_ (.A1(_0569_),
    .A2(_0573_),
    .B1(_0574_),
    .B2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1216_ (.I(_0481_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1217_ (.A1(_0364_),
    .A2(_0362_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1218_ (.I(_0466_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1219_ (.A1(_0582_),
    .A2(_0421_),
    .B1(_0583_),
    .B2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1220_ (.I(_0426_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1221_ (.A1(_0490_),
    .A2(_0585_),
    .B(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1222_ (.I(_0325_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1223_ (.A1(_0264_),
    .A2(_0407_),
    .B(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1224_ (.A1(_0298_),
    .A2(_0258_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1225_ (.A1(_0407_),
    .A2(_0590_),
    .B(_0366_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1226_ (.A1(_0465_),
    .A2(_0389_),
    .A3(_0589_),
    .B1(_0591_),
    .B2(_0475_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1227_ (.I(_0401_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1228_ (.A1(_0570_),
    .A2(_0592_),
    .B(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1229_ (.A1(_0587_),
    .A2(_0592_),
    .B(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1230_ (.A1(_0438_),
    .A2(_0583_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1231_ (.A1(_0267_),
    .A2(_0364_),
    .A3(_0304_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1232_ (.A1(_0584_),
    .A2(_0597_),
    .B(_0472_),
    .C(_0489_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1233_ (.I(_0292_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1234_ (.A1(_0599_),
    .A2(_0385_),
    .B(_0336_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1235_ (.A1(_0363_),
    .A2(_0375_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1236_ (.A1(_0410_),
    .A2(_0521_),
    .B(_0463_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1237_ (.A1(_0280_),
    .A2(_0314_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1238_ (.A1(_0441_),
    .A2(_0557_),
    .B(_0599_),
    .C(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1239_ (.A1(_0601_),
    .A2(_0602_),
    .A3(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1240_ (.A1(_0385_),
    .A2(_0387_),
    .B(_0329_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1241_ (.A1(_0596_),
    .A2(_0598_),
    .A3(_0600_),
    .B1(_0605_),
    .B2(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1242_ (.I(_0455_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1243_ (.A1(_0419_),
    .A2(_0607_),
    .B(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1244_ (.I(_0409_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1245_ (.A1(_0398_),
    .A2(_0582_),
    .B(_0518_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1246_ (.A1(_0255_),
    .A2(_0308_),
    .A3(_0610_),
    .A4(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1247_ (.A1(_0518_),
    .A2(_0522_),
    .B(_0602_),
    .C(_0597_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1248_ (.A1(_0262_),
    .A2(_0289_),
    .A3(_0317_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1249_ (.A1(_0520_),
    .A2(_0508_),
    .A3(_0614_),
    .B(_0292_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1250_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1251_ (.I(_0417_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1252_ (.A1(_0395_),
    .A2(_0616_),
    .B(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1253_ (.A1(_0613_),
    .A2(_0618_),
    .B(_0446_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1254_ (.A1(_0612_),
    .A2(_0619_),
    .B(_0274_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1255_ (.A1(_0595_),
    .A2(_0609_),
    .B(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1256_ (.A1(_0461_),
    .A2(_0555_),
    .B1(_0517_),
    .B2(_0581_),
    .C(_0621_),
    .ZN(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1257_ (.I(_0393_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1258_ (.I(_0369_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1259_ (.A1(_0499_),
    .A2(_0385_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1260_ (.A1(_0623_),
    .A2(_0389_),
    .A3(_0471_),
    .B1(_0624_),
    .B2(_0432_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1261_ (.A1(_0386_),
    .A2(_0324_),
    .A3(_0317_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1262_ (.A1(_0626_),
    .A2(_0375_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1263_ (.A1(_0489_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1264_ (.A1(_0339_),
    .A2(_0320_),
    .B(_0359_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1265_ (.A1(_0528_),
    .A2(_0600_),
    .A3(_0628_),
    .A4(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1266_ (.A1(_0622_),
    .A2(_0625_),
    .B(_0630_),
    .C(_0402_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1267_ (.A1(_0479_),
    .A2(_0280_),
    .A3(_0481_),
    .B(_0527_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1268_ (.A1(_0363_),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1269_ (.A1(_0623_),
    .A2(_0327_),
    .B(_0452_),
    .C(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1270_ (.A1(_0533_),
    .A2(_0388_),
    .A3(_0556_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1271_ (.A1(_0307_),
    .A2(_0519_),
    .B(_0523_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1272_ (.A1(_0424_),
    .A2(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1273_ (.A1(_0540_),
    .A2(_0634_),
    .A3(_0635_),
    .A4(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1274_ (.A1(_0514_),
    .A2(_0631_),
    .A3(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1275_ (.A1(_0535_),
    .A2(_0506_),
    .B(_0293_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1276_ (.A1(_0395_),
    .A2(_0616_),
    .A3(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1277_ (.A1(_0566_),
    .A2(_0434_),
    .A3(_0440_),
    .A4(_0606_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1278_ (.A1(_0333_),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1279_ (.A1(_0544_),
    .A2(_0617_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1280_ (.A1(_0294_),
    .A2(_0320_),
    .A3(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1281_ (.A1(_0641_),
    .A2(_0643_),
    .B(_0645_),
    .C(_0608_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1282_ (.I(_0626_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1283_ (.A1(_0449_),
    .A2(_0293_),
    .A3(_0370_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1284_ (.A1(_0278_),
    .A2(_0488_),
    .B(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1285_ (.A1(_0647_),
    .A2(_0531_),
    .B1(_0649_),
    .B2(_0544_),
    .C(_0501_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1286_ (.A1(_0329_),
    .A2(_0647_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1287_ (.A1(_0315_),
    .A2(_0424_),
    .B1(_0651_),
    .B2(_0442_),
    .C(_0332_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1288_ (.A1(_0537_),
    .A2(_0563_),
    .B(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1289_ (.A1(_0254_),
    .A2(_0479_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1290_ (.A1(_0654_),
    .A2(_0535_),
    .B(_0366_),
    .C(_0599_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1291_ (.A1(_0297_),
    .A2(_0557_),
    .A3(_0278_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1292_ (.A1(_0544_),
    .A2(_0488_),
    .A3(_0655_),
    .A4(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1293_ (.I(_0277_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1294_ (.A1(_0658_),
    .A2(_0288_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1295_ (.A1(_0373_),
    .A2(_0509_),
    .A3(_0614_),
    .B(_0599_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1296_ (.A1(_0399_),
    .A2(_0659_),
    .A3(_0660_),
    .A4(_0651_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1297_ (.A1(_0657_),
    .A2(_0661_),
    .B(_0593_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1298_ (.A1(_0588_),
    .A2(_0494_),
    .B(_0307_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1299_ (.A1(_0312_),
    .A2(_0561_),
    .B1(_0663_),
    .B2(_0534_),
    .C(_0617_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1300_ (.A1(_0335_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1301_ (.A1(_0405_),
    .A2(_0650_),
    .A3(_0653_),
    .B1(_0662_),
    .B2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1302_ (.A1(_0415_),
    .A2(_0454_),
    .B1(_0458_),
    .B2(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1303_ (.A1(_0275_),
    .A2(_0639_),
    .A3(_0646_),
    .B(_0667_),
    .ZN(net10));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1304_ (.A1(_0480_),
    .A2(_0339_),
    .B(_0387_),
    .C(_0658_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1305_ (.A1(_0478_),
    .A2(_0471_),
    .B(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1306_ (.A1(_0495_),
    .A2(_0488_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1307_ (.A1(_0426_),
    .A2(_0603_),
    .A3(_0509_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1308_ (.A1(_0330_),
    .A2(_0670_),
    .B1(_0671_),
    .B2(_0312_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1309_ (.A1(_0452_),
    .A2(_0669_),
    .B(_0672_),
    .C(_0333_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1310_ (.I(_0473_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1311_ (.A1(_0674_),
    .A2(_0378_),
    .A3(_0501_),
    .A4(_0647_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1312_ (.A1(_0525_),
    .A2(_0373_),
    .B(_0577_),
    .C(_0540_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1313_ (.A1(_0405_),
    .A2(_0675_),
    .A3(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1314_ (.A1(_0418_),
    .A2(_0404_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1315_ (.A1(_0437_),
    .A2(_0420_),
    .B1(_0551_),
    .B2(_0406_),
    .C(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1316_ (.A1(_0380_),
    .A2(_0404_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1317_ (.A1(_0453_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1318_ (.A1(_0673_),
    .A2(_0677_),
    .B(_0679_),
    .C(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1319_ (.I(_0445_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1320_ (.A1(_0255_),
    .A2(_0432_),
    .B(_0647_),
    .C(_0674_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1321_ (.A1(_0588_),
    .A2(_0295_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1322_ (.A1(_0555_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1323_ (.A1(_0654_),
    .A2(_0535_),
    .B(_0588_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1324_ (.A1(_0523_),
    .A2(_0687_),
    .B(_0560_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1325_ (.A1(_0302_),
    .A2(_0549_),
    .A3(_0596_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1326_ (.A1(_0399_),
    .A2(_0601_),
    .A3(_0616_),
    .A4(_0640_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1327_ (.A1(_0688_),
    .A2(_0689_),
    .B(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1328_ (.A1(_0644_),
    .A2(_0684_),
    .A3(_0686_),
    .B1(_0691_),
    .B2(_0419_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1329_ (.A1(_0674_),
    .A2(_0437_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1330_ (.A1(_0605_),
    .A2(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1331_ (.A1(_0582_),
    .A2(_0264_),
    .B(_0548_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1332_ (.A1(_0586_),
    .A2(_0596_),
    .A3(_0598_),
    .A4(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1333_ (.A1(_0694_),
    .A2(_0696_),
    .B(_0678_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1334_ (.A1(_0442_),
    .A2(_0526_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1335_ (.A1(_0531_),
    .A2(_0636_),
    .B(_0698_),
    .C(_0550_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1336_ (.A1(_0587_),
    .A2(_0699_),
    .B(_0274_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1337_ (.A1(_0683_),
    .A2(_0692_),
    .B(_0697_),
    .C(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1338_ (.A1(_0461_),
    .A2(_0568_),
    .B1(_0517_),
    .B2(_0682_),
    .C(_0701_),
    .ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1339_ (.A1(_0527_),
    .A2(_0583_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1340_ (.A1(_0685_),
    .A2(_0702_),
    .B(_0566_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1341_ (.A1(_0420_),
    .A2(_0551_),
    .B(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1342_ (.A1(_0449_),
    .A2(_0468_),
    .A3(_0427_),
    .A4(_0451_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1343_ (.A1(_0570_),
    .A2(_0593_),
    .A3(_0648_),
    .B(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1344_ (.A1(_0419_),
    .A2(_0704_),
    .B(_0706_),
    .C(_0273_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1345_ (.A1(_0430_),
    .A2(_0472_),
    .B(_0473_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1346_ (.A1(_0597_),
    .A2(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1347_ (.A1(_0560_),
    .A2(_0495_),
    .A3(_0483_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1348_ (.A1(_0709_),
    .A2(_0710_),
    .B(_0586_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1349_ (.A1(_0482_),
    .A2(_0421_),
    .B(_0648_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1350_ (.A1(_0464_),
    .A2(_0490_),
    .A3(_0712_),
    .B(_0540_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1351_ (.A1(_0278_),
    .A2(_0497_),
    .B(_0498_),
    .C(_0523_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1352_ (.A1(_0407_),
    .A2(_0387_),
    .A3(_0577_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1353_ (.A1(_0494_),
    .A2(_0352_),
    .B(_0714_),
    .C(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1354_ (.A1(_0711_),
    .A2(_0713_),
    .B1(_0716_),
    .B2(_0492_),
    .C(_0273_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1355_ (.A1(_0460_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1356_ (.A1(_0674_),
    .A2(_0522_),
    .A3(_0497_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1357_ (.A1(_0489_),
    .A2(_0474_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1358_ (.A1(_0584_),
    .A2(_0720_),
    .B(_0418_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1359_ (.A1(_0654_),
    .A2(_0421_),
    .A3(_0365_),
    .B1(_0627_),
    .B2(_0623_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1360_ (.A1(_0719_),
    .A2(_0721_),
    .B1(_0722_),
    .B2(_0610_),
    .C(_0427_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1361_ (.A1(_0255_),
    .A2(_0623_),
    .A3(_0432_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1362_ (.A1(_0570_),
    .A2(_0616_),
    .A3(_0640_),
    .A4(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1363_ (.A1(_0723_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1364_ (.A1(_0462_),
    .A2(_0391_),
    .A3(_0357_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1365_ (.A1(_0452_),
    .A2(_0526_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1366_ (.A1(_0302_),
    .A2(_0615_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1367_ (.A1(_0330_),
    .A2(_0670_),
    .B(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1368_ (.A1(_0727_),
    .A2(_0728_),
    .B(_0730_),
    .C(_0333_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1369_ (.A1(_0495_),
    .A2(_0561_),
    .B(_0518_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1370_ (.A1(_0406_),
    .A2(_0429_),
    .B(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1371_ (.A1(_0644_),
    .A2(_0733_),
    .B(_0458_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1372_ (.A1(_0275_),
    .A2(_0726_),
    .B1(_0731_),
    .B2(_0734_),
    .C(_0514_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1373_ (.A1(_0514_),
    .A2(_0707_),
    .A3(_0718_),
    .B(_0735_),
    .ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1374_ (.A1(_0335_),
    .A2(_0675_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1375_ (.A1(_0349_),
    .A2(_0430_),
    .A3(_0374_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1376_ (.A1(_0295_),
    .A2(_0439_),
    .B(_0533_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1377_ (.A1(_0470_),
    .A2(_0370_),
    .B(_0433_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1378_ (.A1(_0439_),
    .A2(_0564_),
    .B1(_0739_),
    .B2(_0327_),
    .C(_0336_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1379_ (.A1(_0566_),
    .A2(_0737_),
    .B(_0738_),
    .C(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1380_ (.A1(_0402_),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1381_ (.A1(_0330_),
    .A2(_0429_),
    .B(_0440_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1382_ (.A1(_0545_),
    .A2(_0743_),
    .B(_0644_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1383_ (.A1(_0736_),
    .A2(_0742_),
    .A3(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1384_ (.A1(_0582_),
    .A2(_0469_),
    .B(_0424_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1385_ (.A1(_0586_),
    .A2(_0649_),
    .B1(_0746_),
    .B2(_0398_),
    .C(_0593_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1386_ (.A1(_0608_),
    .A2(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1387_ (.A1(_0406_),
    .A2(_0521_),
    .B(_0685_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1388_ (.A1(_0622_),
    .A2(_0749_),
    .B(_0680_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1389_ (.A1(_0458_),
    .A2(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1390_ (.A1(_0560_),
    .A2(_0367_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1391_ (.A1(_0353_),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1392_ (.A1(_0371_),
    .A2(_0504_),
    .B1(_0708_),
    .B2(_0327_),
    .C(_0379_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1393_ (.A1(_0629_),
    .A2(_0753_),
    .B1(_0754_),
    .B2(_0610_),
    .C(_0446_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1394_ (.A1(_0480_),
    .A2(_0300_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1395_ (.A1(_0305_),
    .A2(_0408_),
    .B(_0658_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1396_ (.A1(_0409_),
    .A2(_0411_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1397_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1398_ (.A1(_0470_),
    .A2(_0320_),
    .B1(_0507_),
    .B2(_0258_),
    .C(_0527_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1399_ (.A1(_0658_),
    .A2(_0760_),
    .B(_0737_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1400_ (.A1(_0584_),
    .A2(_0597_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1401_ (.A1(_0499_),
    .A2(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1402_ (.A1(_0284_),
    .A2(_0451_),
    .B(_0368_),
    .C(_0336_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1403_ (.A1(_0378_),
    .A2(_0761_),
    .B1(_0763_),
    .B2(_0764_),
    .C(_0617_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1404_ (.A1(_0759_),
    .A2(_0765_),
    .B(_0404_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1405_ (.A1(_0440_),
    .A2(_0606_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1406_ (.A1(_0264_),
    .A2(_0271_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1407_ (.A1(_0480_),
    .A2(_0768_),
    .B1(_0533_),
    .B2(_0321_),
    .C(_0368_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1408_ (.A1(_0303_),
    .A2(_0767_),
    .B(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1409_ (.A1(_0678_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1410_ (.A1(_0460_),
    .A2(_0755_),
    .A3(_0766_),
    .A4(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1411_ (.A1(_0745_),
    .A2(_0748_),
    .A3(_0751_),
    .B1(_0772_),
    .B2(_0516_),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1412_ (.A1(_0610_),
    .A2(_0702_),
    .B(_0683_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1413_ (.A1(_0492_),
    .A2(_0531_),
    .A3(_0474_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1414_ (.A1(_0608_),
    .A2(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1415_ (.I(net3),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1416_ (.A1(_0517_),
    .A2(_0773_),
    .A3(_0775_),
    .B1(_0776_),
    .B2(_0461_),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1417_ (.A1(_0256_),
    .A2(_0314_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1418_ (.I(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1419_ (.I(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1420_ (.I(_0777_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1421_ (.A1(\mod.buffer[134] ),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1422_ (.A1(_0462_),
    .A2(_0779_),
    .B(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1423_ (.I(net1),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1424_ (.I(net6),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1425_ (.A1(_0783_),
    .A2(_0778_),
    .B(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1426_ (.I(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1427_ (.I0(\mod.buffer[133] ),
    .I1(_0782_),
    .S(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1428_ (.I(_0787_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1429_ (.I(_0778_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1430_ (.A1(\mod.buffer[135] ),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1431_ (.A1(_0555_),
    .A2(_0779_),
    .B(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1432_ (.I0(\mod.buffer[134] ),
    .I1(_0790_),
    .S(_0786_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1433_ (.I(_0791_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1434_ (.A1(\mod.buffer[136] ),
    .A2(_0788_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1435_ (.A1(_0622_),
    .A2(_0779_),
    .B(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1436_ (.I(_0785_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1437_ (.I0(\mod.buffer[135] ),
    .I1(_0793_),
    .S(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1438_ (.I(_0795_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1439_ (.A1(\mod.buffer[137] ),
    .A2(_0788_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1440_ (.A1(_0568_),
    .A2(_0780_),
    .B(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1441_ (.I0(\mod.buffer[136] ),
    .I1(_0797_),
    .S(_0794_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1442_ (.I(_0798_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1443_ (.A1(\mod.buffer[138] ),
    .A2(_0788_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1444_ (.A1(_0683_),
    .A2(_0780_),
    .B(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1445_ (.I0(\mod.buffer[137] ),
    .I1(_0800_),
    .S(_0794_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1446_ (.I(_0801_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1447_ (.A1(\mod.buffer[139] ),
    .A2(_0778_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1448_ (.A1(_0516_),
    .A2(_0780_),
    .B(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1449_ (.I0(\mod.buffer[138] ),
    .I1(_0803_),
    .S(_0794_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1450_ (.I(_0804_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1451_ (.A1(_0460_),
    .A2(_0314_),
    .B1(_0779_),
    .B2(net2),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1452_ (.A1(\mod.buffer[139] ),
    .A2(_0786_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1453_ (.A1(_0786_),
    .A2(_0805_),
    .B(_0806_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1454_ (.A1(net6),
    .A2(_0777_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1455_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1456_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1457_ (.I(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1458_ (.I(_0809_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1459_ (.A1(\mod.buffer[7] ),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1460_ (.A1(_0462_),
    .A2(_0810_),
    .B(_0812_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1461_ (.I(_0808_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1462_ (.A1(\mod.buffer[8] ),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1463_ (.A1(_0555_),
    .A2(_0810_),
    .B(_0814_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1464_ (.A1(\mod.buffer[9] ),
    .A2(_0813_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1465_ (.A1(_0622_),
    .A2(_0810_),
    .B(_0815_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1466_ (.A1(\mod.buffer[10] ),
    .A2(_0813_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1467_ (.A1(_0568_),
    .A2(_0810_),
    .B(_0816_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1468_ (.A1(\mod.buffer[11] ),
    .A2(_0813_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1469_ (.A1(_0683_),
    .A2(_0811_),
    .B(_0817_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1470_ (.I(_0808_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1471_ (.A1(\mod.buffer[12] ),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1472_ (.A1(_0516_),
    .A2(_0811_),
    .B(_0819_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1473_ (.A1(\mod.buffer[13] ),
    .A2(_0818_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1474_ (.A1(_0415_),
    .A2(_0811_),
    .B(_0820_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1475_ (.I0(\mod.buffer[7] ),
    .I1(\mod.buffer[14] ),
    .S(_0818_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1476_ (.I(_0821_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1477_ (.I0(\mod.buffer[8] ),
    .I1(\mod.buffer[15] ),
    .S(_0818_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1478_ (.I(_0822_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1479_ (.I(_0809_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1480_ (.I0(\mod.buffer[9] ),
    .I1(\mod.buffer[16] ),
    .S(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1481_ (.I(_0824_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1482_ (.I0(\mod.buffer[10] ),
    .I1(\mod.buffer[17] ),
    .S(_0823_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1483_ (.I(_0825_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1484_ (.I0(\mod.buffer[11] ),
    .I1(\mod.buffer[18] ),
    .S(_0823_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1485_ (.I(_0826_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1486_ (.I0(\mod.buffer[12] ),
    .I1(\mod.buffer[19] ),
    .S(_0823_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1487_ (.I(_0827_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1488_ (.I(_0809_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1489_ (.I0(\mod.buffer[13] ),
    .I1(\mod.buffer[20] ),
    .S(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1490_ (.I(_0829_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1491_ (.I0(\mod.buffer[14] ),
    .I1(\mod.buffer[21] ),
    .S(_0828_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1492_ (.I(_0830_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1493_ (.I0(\mod.buffer[15] ),
    .I1(\mod.buffer[22] ),
    .S(_0828_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1494_ (.I(_0831_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1495_ (.I0(\mod.buffer[16] ),
    .I1(\mod.buffer[23] ),
    .S(_0828_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1496_ (.I(_0832_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1497_ (.I(_0807_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1498_ (.I(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1499_ (.I(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1500_ (.I(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1501_ (.I0(\mod.buffer[17] ),
    .I1(\mod.buffer[24] ),
    .S(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1502_ (.I(_0837_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1503_ (.I0(\mod.buffer[18] ),
    .I1(\mod.buffer[25] ),
    .S(_0836_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1504_ (.I(_0838_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1505_ (.I0(\mod.buffer[19] ),
    .I1(\mod.buffer[26] ),
    .S(_0836_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1506_ (.I(_0839_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1507_ (.I0(\mod.buffer[20] ),
    .I1(\mod.buffer[27] ),
    .S(_0836_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1508_ (.I(_0840_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1509_ (.I(_0835_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1510_ (.I0(\mod.buffer[21] ),
    .I1(\mod.buffer[28] ),
    .S(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1511_ (.I(_0842_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1512_ (.I0(\mod.buffer[22] ),
    .I1(\mod.buffer[29] ),
    .S(_0841_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1513_ (.I(_0843_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1514_ (.I0(\mod.buffer[23] ),
    .I1(\mod.buffer[30] ),
    .S(_0841_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1515_ (.I(_0844_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1516_ (.I0(\mod.buffer[24] ),
    .I1(\mod.buffer[31] ),
    .S(_0841_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1517_ (.I(_0845_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1518_ (.I(_0835_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1519_ (.I0(\mod.buffer[25] ),
    .I1(\mod.buffer[32] ),
    .S(_0846_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1520_ (.I(_0847_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1521_ (.I0(\mod.buffer[26] ),
    .I1(\mod.buffer[33] ),
    .S(_0846_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1522_ (.I(_0848_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1523_ (.I0(\mod.buffer[27] ),
    .I1(\mod.buffer[34] ),
    .S(_0846_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1524_ (.I(_0849_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1525_ (.I0(\mod.buffer[28] ),
    .I1(\mod.buffer[35] ),
    .S(_0846_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1526_ (.I(_0850_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1527_ (.I(_0835_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1528_ (.I0(\mod.buffer[29] ),
    .I1(\mod.buffer[36] ),
    .S(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1529_ (.I(_0852_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1530_ (.I0(\mod.buffer[30] ),
    .I1(\mod.buffer[37] ),
    .S(_0851_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1531_ (.I(_0853_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1532_ (.I0(\mod.buffer[31] ),
    .I1(\mod.buffer[38] ),
    .S(_0851_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1533_ (.I(_0854_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1534_ (.I0(\mod.buffer[32] ),
    .I1(\mod.buffer[39] ),
    .S(_0851_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1535_ (.I(_0855_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1536_ (.I(_0834_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1537_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1538_ (.I0(\mod.buffer[33] ),
    .I1(\mod.buffer[40] ),
    .S(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1539_ (.I(_0858_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1540_ (.I0(\mod.buffer[34] ),
    .I1(\mod.buffer[41] ),
    .S(_0857_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1541_ (.I(_0859_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1542_ (.I0(\mod.buffer[35] ),
    .I1(\mod.buffer[42] ),
    .S(_0857_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1543_ (.I(_0860_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1544_ (.I0(\mod.buffer[36] ),
    .I1(\mod.buffer[43] ),
    .S(_0857_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1545_ (.I(_0861_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1546_ (.I(_0856_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1547_ (.I0(\mod.buffer[37] ),
    .I1(\mod.buffer[44] ),
    .S(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1548_ (.I(_0863_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1549_ (.I0(\mod.buffer[38] ),
    .I1(\mod.buffer[45] ),
    .S(_0862_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1550_ (.I(_0864_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1551_ (.I0(\mod.buffer[39] ),
    .I1(\mod.buffer[46] ),
    .S(_0862_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1552_ (.I(_0865_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1553_ (.I0(\mod.buffer[40] ),
    .I1(\mod.buffer[47] ),
    .S(_0862_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1554_ (.I(_0866_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1555_ (.I(_0856_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1556_ (.I0(\mod.buffer[41] ),
    .I1(\mod.buffer[48] ),
    .S(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1557_ (.I(_0868_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1558_ (.I0(\mod.buffer[42] ),
    .I1(\mod.buffer[49] ),
    .S(_0867_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1559_ (.I(_0869_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1560_ (.I0(\mod.buffer[43] ),
    .I1(\mod.buffer[50] ),
    .S(_0867_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1561_ (.I(_0870_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1562_ (.I0(\mod.buffer[44] ),
    .I1(\mod.buffer[51] ),
    .S(_0867_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1563_ (.I(_0871_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1564_ (.I(_0856_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1565_ (.I0(\mod.buffer[45] ),
    .I1(\mod.buffer[52] ),
    .S(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1566_ (.I(_0873_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1567_ (.I0(\mod.buffer[46] ),
    .I1(\mod.buffer[53] ),
    .S(_0872_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1568_ (.I(_0874_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1569_ (.I0(\mod.buffer[47] ),
    .I1(\mod.buffer[54] ),
    .S(_0872_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1570_ (.I(_0875_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1571_ (.I0(\mod.buffer[48] ),
    .I1(\mod.buffer[55] ),
    .S(_0872_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1572_ (.I(_0876_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1573_ (.I(_0834_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1574_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1575_ (.I0(\mod.buffer[49] ),
    .I1(\mod.buffer[56] ),
    .S(_0878_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1576_ (.I(_0879_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1577_ (.I0(\mod.buffer[50] ),
    .I1(\mod.buffer[57] ),
    .S(_0878_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1578_ (.I(_0880_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1579_ (.I0(\mod.buffer[51] ),
    .I1(\mod.buffer[58] ),
    .S(_0878_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1580_ (.I(_0146_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1581_ (.I0(\mod.buffer[52] ),
    .I1(\mod.buffer[59] ),
    .S(_0878_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1582_ (.I(_0147_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1583_ (.I(_0877_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1584_ (.I0(\mod.buffer[53] ),
    .I1(\mod.buffer[60] ),
    .S(_0148_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1585_ (.I(_0149_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1586_ (.I0(\mod.buffer[54] ),
    .I1(\mod.buffer[61] ),
    .S(_0148_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1587_ (.I(_0150_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1588_ (.I0(\mod.buffer[55] ),
    .I1(\mod.buffer[62] ),
    .S(_0148_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1589_ (.I(_0151_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1590_ (.I0(\mod.buffer[56] ),
    .I1(\mod.buffer[63] ),
    .S(_0148_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1591_ (.I(_0152_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1592_ (.I(_0877_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1593_ (.I0(\mod.buffer[57] ),
    .I1(\mod.buffer[64] ),
    .S(_0153_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1594_ (.I(_0154_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1595_ (.I0(\mod.buffer[58] ),
    .I1(\mod.buffer[65] ),
    .S(_0153_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1596_ (.I(_0155_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1597_ (.I0(\mod.buffer[59] ),
    .I1(\mod.buffer[66] ),
    .S(_0153_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1598_ (.I(_0156_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1599_ (.I0(\mod.buffer[60] ),
    .I1(\mod.buffer[67] ),
    .S(_0153_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1600_ (.I(_0157_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1601_ (.I(_0877_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1602_ (.I0(\mod.buffer[61] ),
    .I1(\mod.buffer[68] ),
    .S(_0158_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1603_ (.I(_0159_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1604_ (.I0(\mod.buffer[62] ),
    .I1(\mod.buffer[69] ),
    .S(_0158_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1605_ (.I(_0160_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1606_ (.I0(\mod.buffer[63] ),
    .I1(\mod.buffer[70] ),
    .S(_0158_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1607_ (.I(_0161_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1608_ (.I0(\mod.buffer[64] ),
    .I1(\mod.buffer[71] ),
    .S(_0158_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1609_ (.I(_0162_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1610_ (.I(_0834_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1611_ (.I(_0163_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1612_ (.I0(\mod.buffer[65] ),
    .I1(\mod.buffer[72] ),
    .S(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1613_ (.I(_0165_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1614_ (.I0(\mod.buffer[66] ),
    .I1(\mod.buffer[73] ),
    .S(_0164_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1615_ (.I(_0166_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1616_ (.I0(\mod.buffer[67] ),
    .I1(\mod.buffer[74] ),
    .S(_0164_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1617_ (.I(_0167_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1618_ (.I0(\mod.buffer[68] ),
    .I1(\mod.buffer[75] ),
    .S(_0164_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1619_ (.I(_0168_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1620_ (.I(_0163_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1621_ (.I0(\mod.buffer[69] ),
    .I1(\mod.buffer[76] ),
    .S(_0169_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1622_ (.I(_0170_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1623_ (.I0(\mod.buffer[70] ),
    .I1(\mod.buffer[77] ),
    .S(_0169_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1624_ (.I(_0171_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1625_ (.I0(\mod.buffer[71] ),
    .I1(\mod.buffer[78] ),
    .S(_0169_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1626_ (.I(_0172_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1627_ (.I0(\mod.buffer[72] ),
    .I1(\mod.buffer[79] ),
    .S(_0169_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1628_ (.I(_0173_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1629_ (.I(_0163_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1630_ (.I0(\mod.buffer[73] ),
    .I1(\mod.buffer[80] ),
    .S(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1631_ (.I(_0175_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1632_ (.I0(\mod.buffer[74] ),
    .I1(\mod.buffer[81] ),
    .S(_0174_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1633_ (.I(_0176_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1634_ (.I0(\mod.buffer[75] ),
    .I1(\mod.buffer[82] ),
    .S(_0174_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1635_ (.I(_0177_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1636_ (.I0(\mod.buffer[76] ),
    .I1(\mod.buffer[83] ),
    .S(_0174_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1637_ (.I(_0178_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1638_ (.I(_0163_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1639_ (.I0(\mod.buffer[77] ),
    .I1(\mod.buffer[84] ),
    .S(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1640_ (.I(_0180_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1641_ (.I0(\mod.buffer[78] ),
    .I1(\mod.buffer[85] ),
    .S(_0179_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1642_ (.I(_0181_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1643_ (.I0(\mod.buffer[79] ),
    .I1(\mod.buffer[86] ),
    .S(_0179_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1644_ (.I(_0182_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1645_ (.I0(\mod.buffer[80] ),
    .I1(\mod.buffer[87] ),
    .S(_0179_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1646_ (.I(_0183_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1647_ (.I(_0833_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1648_ (.I(_0184_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1649_ (.I0(\mod.buffer[81] ),
    .I1(\mod.buffer[88] ),
    .S(_0185_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1650_ (.I(_0186_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1651_ (.I0(\mod.buffer[82] ),
    .I1(\mod.buffer[89] ),
    .S(_0185_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1652_ (.I(_0187_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1653_ (.I0(\mod.buffer[83] ),
    .I1(\mod.buffer[90] ),
    .S(_0185_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1654_ (.I(_0188_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1655_ (.I0(\mod.buffer[84] ),
    .I1(\mod.buffer[91] ),
    .S(_0185_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1656_ (.I(_0189_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1657_ (.I(_0184_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1658_ (.I0(\mod.buffer[85] ),
    .I1(\mod.buffer[92] ),
    .S(_0190_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1659_ (.I(_0191_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1660_ (.I0(\mod.buffer[86] ),
    .I1(\mod.buffer[93] ),
    .S(_0190_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1661_ (.I(_0192_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1662_ (.I0(\mod.buffer[87] ),
    .I1(\mod.buffer[94] ),
    .S(_0190_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1663_ (.I(_0193_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1664_ (.I0(\mod.buffer[88] ),
    .I1(\mod.buffer[95] ),
    .S(_0190_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1665_ (.I(_0194_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1666_ (.I(_0184_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1667_ (.I0(\mod.buffer[89] ),
    .I1(\mod.buffer[96] ),
    .S(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1668_ (.I(_0196_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1669_ (.I0(\mod.buffer[90] ),
    .I1(\mod.buffer[97] ),
    .S(_0195_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1670_ (.I(_0197_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1671_ (.I0(\mod.buffer[91] ),
    .I1(\mod.buffer[98] ),
    .S(_0195_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1672_ (.I(_0198_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1673_ (.I0(\mod.buffer[92] ),
    .I1(\mod.buffer[99] ),
    .S(_0195_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1674_ (.I(_0199_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1675_ (.I(_0184_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1676_ (.I0(\mod.buffer[93] ),
    .I1(\mod.buffer[100] ),
    .S(_0200_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1677_ (.I(_0201_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1678_ (.I0(\mod.buffer[94] ),
    .I1(\mod.buffer[101] ),
    .S(_0200_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1679_ (.I(_0202_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1680_ (.I0(\mod.buffer[95] ),
    .I1(\mod.buffer[102] ),
    .S(_0200_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1681_ (.I(_0203_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1682_ (.I0(\mod.buffer[96] ),
    .I1(\mod.buffer[103] ),
    .S(_0200_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1683_ (.I(_0204_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1684_ (.I(_0833_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1685_ (.I(_0205_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1686_ (.I0(\mod.buffer[97] ),
    .I1(\mod.buffer[104] ),
    .S(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1687_ (.I(_0207_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1688_ (.I0(\mod.buffer[98] ),
    .I1(\mod.buffer[105] ),
    .S(_0206_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1689_ (.I(_0208_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1690_ (.I0(\mod.buffer[99] ),
    .I1(\mod.buffer[106] ),
    .S(_0206_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1691_ (.I(_0209_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1692_ (.I0(\mod.buffer[100] ),
    .I1(\mod.buffer[107] ),
    .S(_0206_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1693_ (.I(_0210_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1694_ (.I(_0205_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1695_ (.I0(\mod.buffer[101] ),
    .I1(\mod.buffer[108] ),
    .S(_0211_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1696_ (.I(_0212_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1697_ (.I0(\mod.buffer[102] ),
    .I1(\mod.buffer[109] ),
    .S(_0211_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1698_ (.I(_0213_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1699_ (.I0(\mod.buffer[103] ),
    .I1(\mod.buffer[110] ),
    .S(_0211_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1700_ (.I(_0214_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1701_ (.I0(\mod.buffer[104] ),
    .I1(\mod.buffer[111] ),
    .S(_0211_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1702_ (.I(_0215_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1703_ (.I(_0205_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1704_ (.I0(\mod.buffer[105] ),
    .I1(\mod.buffer[112] ),
    .S(_0216_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1705_ (.I(_0217_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1706_ (.I0(\mod.buffer[106] ),
    .I1(\mod.buffer[113] ),
    .S(_0216_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1707_ (.I(_0218_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1708_ (.I0(\mod.buffer[107] ),
    .I1(\mod.buffer[114] ),
    .S(_0216_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1709_ (.I(_0219_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1710_ (.I0(\mod.buffer[108] ),
    .I1(\mod.buffer[115] ),
    .S(_0216_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1711_ (.I(_0220_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1712_ (.I(_0205_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1713_ (.I0(\mod.buffer[109] ),
    .I1(\mod.buffer[116] ),
    .S(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1714_ (.I(_0222_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1715_ (.I0(\mod.buffer[110] ),
    .I1(\mod.buffer[117] ),
    .S(_0221_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1716_ (.I(_0223_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1717_ (.I0(\mod.buffer[111] ),
    .I1(\mod.buffer[118] ),
    .S(_0221_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1718_ (.I(_0224_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1719_ (.I0(\mod.buffer[112] ),
    .I1(\mod.buffer[119] ),
    .S(_0221_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1720_ (.I(_0225_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1721_ (.I(_0833_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1722_ (.I(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1723_ (.I0(\mod.buffer[113] ),
    .I1(\mod.buffer[120] ),
    .S(_0227_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1724_ (.I(_0228_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1725_ (.I0(\mod.buffer[114] ),
    .I1(\mod.buffer[121] ),
    .S(_0227_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1726_ (.I(_0229_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1727_ (.I0(\mod.buffer[115] ),
    .I1(\mod.buffer[122] ),
    .S(_0227_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1728_ (.I(_0230_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1729_ (.I0(\mod.buffer[116] ),
    .I1(\mod.buffer[123] ),
    .S(_0227_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1730_ (.I(_0231_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1731_ (.I(_0226_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1732_ (.I0(\mod.buffer[117] ),
    .I1(\mod.buffer[124] ),
    .S(_0232_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1733_ (.I(_0233_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1734_ (.I0(\mod.buffer[118] ),
    .I1(\mod.buffer[125] ),
    .S(_0232_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1735_ (.I(_0234_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1736_ (.I0(\mod.buffer[119] ),
    .I1(\mod.buffer[126] ),
    .S(_0232_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1737_ (.I(_0235_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1738_ (.I0(\mod.buffer[120] ),
    .I1(\mod.buffer[127] ),
    .S(_0232_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1739_ (.I(_0236_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1740_ (.I(_0226_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1741_ (.I0(\mod.buffer[121] ),
    .I1(\mod.buffer[128] ),
    .S(_0237_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1742_ (.I(_0238_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1743_ (.I0(\mod.buffer[122] ),
    .I1(\mod.buffer[129] ),
    .S(_0237_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1744_ (.I(_0239_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1745_ (.I0(\mod.buffer[123] ),
    .I1(\mod.buffer[130] ),
    .S(_0237_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1746_ (.I(_0240_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1747_ (.I0(\mod.buffer[124] ),
    .I1(\mod.buffer[131] ),
    .S(_0237_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1748_ (.I(_0241_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1749_ (.I(_0226_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1750_ (.I0(\mod.buffer[125] ),
    .I1(\mod.buffer[132] ),
    .S(_0242_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1751_ (.I(_0243_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1752_ (.I0(\mod.buffer[126] ),
    .I1(\mod.buffer[133] ),
    .S(_0242_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1753_ (.I(_0244_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1754_ (.I0(\mod.buffer[127] ),
    .I1(\mod.buffer[134] ),
    .S(_0242_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1755_ (.I(_0245_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1756_ (.I0(\mod.buffer[128] ),
    .I1(\mod.buffer[135] ),
    .S(_0242_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1757_ (.I(_0246_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1758_ (.I(_0808_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1759_ (.I0(\mod.buffer[129] ),
    .I1(\mod.buffer[136] ),
    .S(_0247_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1760_ (.I(_0248_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1761_ (.I0(\mod.buffer[130] ),
    .I1(\mod.buffer[137] ),
    .S(_0247_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1762_ (.I(_0249_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1763_ (.I0(\mod.buffer[131] ),
    .I1(\mod.buffer[138] ),
    .S(_0247_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1764_ (.I(_0250_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1765_ (.I0(\mod.buffer[132] ),
    .I1(\mod.buffer[139] ),
    .S(_0247_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1766_ (.I(_0251_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1767_ (.I(_0784_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1768_ (.I(_0784_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1769_ (.I(_0784_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1770_ (.D(_0006_),
    .CLK(net16),
    .Q(\mod.buffer[133] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1771_ (.D(_0007_),
    .CLK(net16),
    .Q(\mod.buffer[134] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1772_ (.D(_0008_),
    .CLK(net17),
    .Q(\mod.buffer[135] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1773_ (.D(_0009_),
    .CLK(net27),
    .Q(\mod.buffer[136] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1774_ (.D(_0010_),
    .CLK(net23),
    .Q(\mod.buffer[137] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1775_ (.D(_0011_),
    .CLK(net27),
    .Q(\mod.buffer[138] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1776_ (.D(_0012_),
    .CLK(net17),
    .Q(\mod.buffer[139] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1777_ (.D(_0013_),
    .CLK(net15),
    .Q(\mod.buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1778_ (.D(_0014_),
    .CLK(net27),
    .Q(\mod.buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1779_ (.D(_0015_),
    .CLK(net48),
    .Q(\mod.buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1780_ (.D(_0016_),
    .CLK(net48),
    .Q(\mod.buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1781_ (.D(_0017_),
    .CLK(net48),
    .Q(\mod.buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1782_ (.D(_0018_),
    .CLK(net47),
    .Q(\mod.buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1783_ (.D(_0019_),
    .CLK(net47),
    .Q(\mod.buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1784_ (.D(_0020_),
    .CLK(net47),
    .Q(\mod.buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1785_ (.D(_0021_),
    .CLK(net43),
    .Q(\mod.buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1786_ (.D(_0022_),
    .CLK(net50),
    .Q(\mod.buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1787_ (.D(_0023_),
    .CLK(net48),
    .Q(\mod.buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1788_ (.D(_0024_),
    .CLK(net49),
    .Q(\mod.buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1789_ (.D(_0025_),
    .CLK(net49),
    .Q(\mod.buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1790_ (.D(_0026_),
    .CLK(net45),
    .Q(\mod.buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1791_ (.D(_0027_),
    .CLK(net43),
    .Q(\mod.buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1792_ (.D(_0028_),
    .CLK(net43),
    .Q(\mod.buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1793_ (.D(_0029_),
    .CLK(net45),
    .Q(\mod.buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1794_ (.D(_0030_),
    .CLK(net49),
    .Q(\mod.buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1795_ (.D(_0031_),
    .CLK(net51),
    .Q(\mod.buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1796_ (.D(_0032_),
    .CLK(net54),
    .Q(\mod.buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1797_ (.D(_0033_),
    .CLK(net50),
    .Q(\mod.buffer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1798_ (.D(_0034_),
    .CLK(net50),
    .Q(\mod.buffer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1799_ (.D(_0035_),
    .CLK(net43),
    .Q(\mod.buffer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1800_ (.D(_0036_),
    .CLK(net45),
    .Q(\mod.buffer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1801_ (.D(_0037_),
    .CLK(net50),
    .Q(\mod.buffer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1802_ (.D(_0038_),
    .CLK(net51),
    .Q(\mod.buffer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1803_ (.D(_0039_),
    .CLK(net51),
    .Q(\mod.buffer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1804_ (.D(_0040_),
    .CLK(net51),
    .Q(\mod.buffer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1805_ (.D(_0041_),
    .CLK(net52),
    .Q(\mod.buffer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1806_ (.D(_0042_),
    .CLK(net44),
    .Q(\mod.buffer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1807_ (.D(_0043_),
    .CLK(net45),
    .Q(\mod.buffer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1808_ (.D(_0044_),
    .CLK(net53),
    .Q(\mod.buffer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1809_ (.D(_0045_),
    .CLK(net52),
    .Q(\mod.buffer[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1810_ (.D(_0046_),
    .CLK(net65),
    .Q(\mod.buffer[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1811_ (.D(_0047_),
    .CLK(net65),
    .Q(\mod.buffer[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1812_ (.D(_0048_),
    .CLK(net52),
    .Q(\mod.buffer[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1813_ (.D(_0049_),
    .CLK(net46),
    .Q(\mod.buffer[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1814_ (.D(_0050_),
    .CLK(net56),
    .Q(\mod.buffer[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1815_ (.D(_0051_),
    .CLK(net64),
    .Q(\mod.buffer[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1816_ (.D(_0052_),
    .CLK(net65),
    .Q(\mod.buffer[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1817_ (.D(_0053_),
    .CLK(net65),
    .Q(\mod.buffer[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1818_ (.D(_0054_),
    .CLK(net66),
    .Q(\mod.buffer[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1819_ (.D(_0055_),
    .CLK(net64),
    .Q(\mod.buffer[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1820_ (.D(_0056_),
    .CLK(net58),
    .Q(\mod.buffer[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1821_ (.D(_0057_),
    .CLK(net56),
    .Q(\mod.buffer[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1822_ (.D(_0058_),
    .CLK(net64),
    .Q(\mod.buffer[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1823_ (.D(_0059_),
    .CLK(net66),
    .Q(\mod.buffer[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1824_ (.D(_0060_),
    .CLK(net70),
    .Q(\mod.buffer[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1825_ (.D(_0061_),
    .CLK(net70),
    .Q(\mod.buffer[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1826_ (.D(_0062_),
    .CLK(net64),
    .Q(\mod.buffer[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1827_ (.D(_0063_),
    .CLK(net58),
    .Q(\mod.buffer[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1828_ (.D(_0064_),
    .CLK(net57),
    .Q(\mod.buffer[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1829_ (.D(_0065_),
    .CLK(net67),
    .Q(\mod.buffer[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1830_ (.D(_0066_),
    .CLK(net68),
    .Q(\mod.buffer[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1831_ (.D(_0067_),
    .CLK(net68),
    .Q(\mod.buffer[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1832_ (.D(_0068_),
    .CLK(net68),
    .Q(\mod.buffer[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1833_ (.D(_0069_),
    .CLK(net69),
    .Q(\mod.buffer[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1834_ (.D(_0070_),
    .CLK(net61),
    .Q(\mod.buffer[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1835_ (.D(_0071_),
    .CLK(net58),
    .Q(\mod.buffer[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1836_ (.D(_0072_),
    .CLK(net63),
    .Q(\mod.buffer[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1837_ (.D(_0073_),
    .CLK(net68),
    .Q(\mod.buffer[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1838_ (.D(_0074_),
    .CLK(net61),
    .Q(\mod.buffer[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1839_ (.D(_0075_),
    .CLK(net69),
    .Q(\mod.buffer[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1840_ (.D(_0076_),
    .CLK(net61),
    .Q(\mod.buffer[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1841_ (.D(_0077_),
    .CLK(net61),
    .Q(\mod.buffer[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1842_ (.D(_0078_),
    .CLK(net59),
    .Q(\mod.buffer[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1843_ (.D(_0079_),
    .CLK(net57),
    .Q(\mod.buffer[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1844_ (.D(_0080_),
    .CLK(net59),
    .Q(\mod.buffer[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1845_ (.D(_0081_),
    .CLK(net62),
    .Q(\mod.buffer[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1846_ (.D(_0082_),
    .CLK(net60),
    .Q(\mod.buffer[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1847_ (.D(_0083_),
    .CLK(net60),
    .Q(\mod.buffer[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1848_ (.D(_0084_),
    .CLK(net60),
    .Q(\mod.buffer[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1849_ (.D(_0085_),
    .CLK(net59),
    .Q(\mod.buffer[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1850_ (.D(_0086_),
    .CLK(net57),
    .Q(\mod.buffer[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1851_ (.D(_0087_),
    .CLK(net59),
    .Q(\mod.buffer[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1852_ (.D(_0088_),
    .CLK(net37),
    .Q(\mod.buffer[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1853_ (.D(_0089_),
    .CLK(net37),
    .Q(\mod.buffer[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1854_ (.D(_0090_),
    .CLK(net38),
    .Q(\mod.buffer[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1855_ (.D(_0091_),
    .CLK(net38),
    .Q(\mod.buffer[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1856_ (.D(_0092_),
    .CLK(net35),
    .Q(\mod.buffer[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1857_ (.D(_0093_),
    .CLK(net33),
    .Q(\mod.buffer[80] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1858_ (.D(_0094_),
    .CLK(net37),
    .Q(\mod.buffer[81] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1859_ (.D(_0095_),
    .CLK(net36),
    .Q(\mod.buffer[82] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1860_ (.D(_0096_),
    .CLK(net36),
    .Q(\mod.buffer[83] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1861_ (.D(_0097_),
    .CLK(net32),
    .Q(\mod.buffer[84] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1862_ (.D(_0098_),
    .CLK(net35),
    .Q(\mod.buffer[85] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1863_ (.D(_0099_),
    .CLK(net33),
    .Q(\mod.buffer[86] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1864_ (.D(_0100_),
    .CLK(net34),
    .Q(\mod.buffer[87] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1865_ (.D(_0101_),
    .CLK(net37),
    .Q(\mod.buffer[88] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1866_ (.D(_0102_),
    .CLK(net35),
    .Q(\mod.buffer[89] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1867_ (.D(_0103_),
    .CLK(net32),
    .Q(\mod.buffer[90] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1868_ (.D(_0104_),
    .CLK(net32),
    .Q(\mod.buffer[91] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1869_ (.D(_0105_),
    .CLK(net35),
    .Q(\mod.buffer[92] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1870_ (.D(_0106_),
    .CLK(net33),
    .Q(\mod.buffer[93] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1871_ (.D(_0107_),
    .CLK(net56),
    .Q(\mod.buffer[94] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1872_ (.D(_0108_),
    .CLK(net34),
    .Q(\mod.buffer[95] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1873_ (.D(_0109_),
    .CLK(net30),
    .Q(\mod.buffer[96] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1874_ (.D(_0110_),
    .CLK(net30),
    .Q(\mod.buffer[97] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1875_ (.D(_0111_),
    .CLK(net30),
    .Q(\mod.buffer[98] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1876_ (.D(_0112_),
    .CLK(net30),
    .Q(\mod.buffer[99] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1877_ (.D(_0113_),
    .CLK(net33),
    .Q(\mod.buffer[100] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1878_ (.D(_0114_),
    .CLK(net56),
    .Q(\mod.buffer[101] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1879_ (.D(_0115_),
    .CLK(net34),
    .Q(\mod.buffer[102] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1880_ (.D(_0116_),
    .CLK(net29),
    .Q(\mod.buffer[103] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1881_ (.D(_0117_),
    .CLK(net31),
    .Q(\mod.buffer[104] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1882_ (.D(_0118_),
    .CLK(net29),
    .Q(\mod.buffer[105] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1883_ (.D(_0119_),
    .CLK(net29),
    .Q(\mod.buffer[106] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1884_ (.D(_0120_),
    .CLK(net23),
    .Q(\mod.buffer[107] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1885_ (.D(_0121_),
    .CLK(net44),
    .Q(\mod.buffer[108] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1886_ (.D(_0122_),
    .CLK(net24),
    .Q(\mod.buffer[109] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1887_ (.D(_0123_),
    .CLK(net29),
    .Q(\mod.buffer[110] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1888_ (.D(_0124_),
    .CLK(net31),
    .Q(\mod.buffer[111] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1889_ (.D(_0125_),
    .CLK(net19),
    .Q(\mod.buffer[112] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1890_ (.D(_0126_),
    .CLK(net20),
    .Q(\mod.buffer[113] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1891_ (.D(_0127_),
    .CLK(net26),
    .Q(\mod.buffer[114] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1892_ (.D(_0128_),
    .CLK(net25),
    .Q(\mod.buffer[115] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1893_ (.D(_0129_),
    .CLK(net25),
    .Q(\mod.buffer[116] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1894_ (.D(_0130_),
    .CLK(net20),
    .Q(\mod.buffer[117] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1895_ (.D(_0131_),
    .CLK(net19),
    .Q(\mod.buffer[118] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1896_ (.D(_0132_),
    .CLK(net21),
    .Q(\mod.buffer[119] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1897_ (.D(_0133_),
    .CLK(net18),
    .Q(\mod.buffer[120] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1898_ (.D(_0134_),
    .CLK(net23),
    .Q(\mod.buffer[121] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1899_ (.D(_0135_),
    .CLK(net24),
    .Q(\mod.buffer[122] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1900_ (.D(_0136_),
    .CLK(net24),
    .Q(\mod.buffer[123] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1901_ (.D(_0137_),
    .CLK(net21),
    .Q(\mod.buffer[124] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1902_ (.D(_0138_),
    .CLK(net18),
    .Q(\mod.buffer[125] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1903_ (.D(_0139_),
    .CLK(net18),
    .Q(\mod.buffer[126] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1904_ (.D(_0140_),
    .CLK(net19),
    .Q(\mod.buffer[127] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1905_ (.D(_0141_),
    .CLK(net20),
    .Q(\mod.buffer[128] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1906_ (.D(_0142_),
    .CLK(net24),
    .Q(\mod.buffer[129] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1907_ (.D(_0143_),
    .CLK(net23),
    .Q(\mod.buffer[130] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1908_ (.D(_0144_),
    .CLK(net20),
    .Q(\mod.buffer[131] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1909_ (.D(_0145_),
    .CLK(net18),
    .Q(\mod.buffer[132] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1910_ (.D(_0000_),
    .RN(_0003_),
    .CLK(net15),
    .Q(\mod.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1911_ (.D(_0001_),
    .RN(_0004_),
    .CLK(net15),
    .Q(\mod.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1912_ (.D(_0002_),
    .RN(_0005_),
    .CLK(net15),
    .Q(\mod.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__D (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[8]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(io_in[9]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output9 (.I(net9),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout15 (.I(net17),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout16 (.I(net17),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout17 (.I(net22),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout18 (.I(net19),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout19 (.I(net21),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout20 (.I(net21),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout21 (.I(net22),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout22 (.I(net28),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout23 (.I(net26),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout24 (.I(net26),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout25 (.I(net26),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout26 (.I(net27),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout27 (.I(net28),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout28 (.I(net42),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout29 (.I(net31),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout32 (.I(net41),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout33 (.I(net40),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout34 (.I(net40),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout35 (.I(net39),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout36 (.I(net39),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout37 (.I(net39),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout38 (.I(net39),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net74),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net46),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net46),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net47),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net55),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net54),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout50 (.I(net53),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net53),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net73),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net63),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout59 (.I(net62),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net62),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net63),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net72),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout64 (.I(net67),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout65 (.I(net67),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net71),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout68 (.I(net70),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net71),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net74),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net5),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__S (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__S (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__S (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__S (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__S (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__S (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__S (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__S (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__S (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__S (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__S (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__S (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__S (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__S (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__S (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__S (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__S (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__S (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__S (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__S (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__S (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__S (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__S (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__S (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__S (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__S (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__S (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__S (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__S (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__S (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__S (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__S (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__S (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__S (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__S (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__S (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__S (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__S (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__S (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__S (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__S (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__S (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__S (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__S (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__S (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__S (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__S (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__S (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__S (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__S (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__S (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__S (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__S (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__S (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__S (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__S (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__S (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__S (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__S (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__S (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1320__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0886__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1417__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__B (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0890__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0886__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__B2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1224__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0889__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1100__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0890__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1140__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0930__I (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A2 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0992__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0895__I (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A1 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1331__A2 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__A1 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__A1 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0938__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0928__I (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0913__I (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0897__I (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1231__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0927__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__I0 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A2 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__A2 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__A2 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__C (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1344__C (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1090__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1336__B (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1254__B (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0907__I (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0994__I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0942__I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0909__I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__A3 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1284__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1267__A2 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1000__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1197__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1070__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0947__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0925__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1249__B (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1233__I (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1065__I (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0925__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1085__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__B1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0932__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1107__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0931__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__B2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__A1 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__A1 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1086__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__C (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1231__A3 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1156__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__B (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0937__I (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1395__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1095__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1298__B (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1271__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__A3 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__B (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1042__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0943__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1308__B2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1299__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__B2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1031__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1417__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0947__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1287__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1069__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1107__A3 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0951__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1000__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A3 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A4 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1107__A2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1073__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1120__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A4 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0958__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__B2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1378__B2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__B (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1286__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1240__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1072__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0962__I (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1381__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1308__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__B2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1287__C (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__C (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1125__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0965__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__C (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__C (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1278__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__C (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1300__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1214__B (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1014__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__C (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1378__C (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__B (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1160__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1153__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0971__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1304__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__A3 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1118__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1019__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__A3 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1131__B (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1074__I (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1058__I (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0984__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1353__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1185__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__B (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1156__A3 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1131__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1127__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1168__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1159__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__C (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1364__A3 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__B (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1038__I (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1231__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1217__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1026__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1390__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__C (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__B (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__A3 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1258__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1198__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1026__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1201__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__B2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1145__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__B3 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1145__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__B2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__C (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__I (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__I (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1316__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__C (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1088__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__C (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1240__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1020__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1304__B (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1240__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1020__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1145__A3 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1026__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1023__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1364__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1192__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1177__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1167__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1027__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1027__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1276__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1144__B (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1035__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1190__B (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1043__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1385__B2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__B2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1296__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__C (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1227__I (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__I (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__C (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__C (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1035__C (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1316__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1314__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1037__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1313__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1136__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1045__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1387__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__B2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1044__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1225__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__I (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1044__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1236__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1159__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1111__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1043__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1045__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1092__A2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__B (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1314__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1183__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1051__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1341__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1359__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A3 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__B (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1287__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A4 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__C (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1068__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1171__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1120__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1084__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1061__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1381__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1085__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1130__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1064__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__B (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1167__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1277__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__A4 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1329__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1071__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1378__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1199__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1072__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1381__B (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1277__A3 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__B1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1199__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__B2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1287__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1129__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__C (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__C (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1253__B (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1079__C (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1130__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__A4 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1084__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1365__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__B (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1302__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1203__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__B2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1242__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1183__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__C (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1088__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1410__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1094__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__B2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1256__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1188__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1364__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1188__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1236__B (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1097__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1124__C (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1110__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__I (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1109__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1190__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1104__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1131__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1104__B (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__A3 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1109__A3 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__B (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__A3 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1109__B1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__B (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1310__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1151__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__A3 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__A1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__A1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1135__A1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1124__A1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1289__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1267__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1304__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1267__A3 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1115__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__B2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1190__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1128__I (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1123__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__C (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1123__B (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1124__B (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__B2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1146__B2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1126__B (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1148__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__A3 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1133__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1401__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1144__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1133__B (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__A3 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__C (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__C (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1135__C (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__A3 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__B (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1148__B1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__C (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1148__B2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1411__B2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1150__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__B1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1256__B1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__B (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1247__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__B (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1271__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1192__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1153__A3 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1387__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1236__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__B (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__A2 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1247__A2 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__A2 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__A3 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__C (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1324__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1271__B (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__A4 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1169__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1159__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1365__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__C (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1267__B (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1161__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__B2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__B1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__B (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1270__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1205__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__B2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1288__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1210__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1171__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__B (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__C (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__B2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1292__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__B2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1279__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__A3 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1331__B (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1341__A2 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__A2 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1185__A2 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1322__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1256__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1192__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1390__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1347__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1324__B (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1196__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1299__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__B1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1196__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1288__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1198__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__B (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1277__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1201__C (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1203__C (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__A3 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__B (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1331__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1245__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__B1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__B2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1336__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1323__B (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1298__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__B (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__B1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1385__C (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1297__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1247__C (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__B (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1290__C (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1238__B (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1265__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__A3 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1277__A4 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__B2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1414__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__C (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1243__B (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__B2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__B2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A3 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__A3 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1249__A3 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1250__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__C (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1299__C (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1279__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__B (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1256__C (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1435__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1388__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1359__B2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__B (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__C (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__A3 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__A3 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__A4 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1276__A3 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1328__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__A3 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1320__B (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__A4 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1286__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__A3 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1284__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1385__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__B1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__A3 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1359__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1323__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1290__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1296__A3 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1308__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1308__B1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1329__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1320__C (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1333__B (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__C (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__B (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1337__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1333__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__B1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__B1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__B (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__B (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__B (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1378__B1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1411__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1411__A3 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1401__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A2 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__B1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1421__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__B (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__S (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__S (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__S (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__S (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1466__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1486__S (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__S (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__S (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__S (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__S (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__S (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__S (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__S (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1499__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__I (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__I (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__I (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__I (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__S (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__S (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__S (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__S (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__S (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__S (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__S (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__S (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__S (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__S (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__S (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__S (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__S (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__S (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__S (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__S (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__S (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__S (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__S (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__S (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__S (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__S (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__S (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__S (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__S (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__S (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__S (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__S (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__S (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1015__I (.I(\mod.buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0956__I (.I(\mod.buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0921__I (.I(\mod.buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__I (.I(\mod.buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__I0 (.I(\mod.buffer[104] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__I1 (.I(\mod.buffer[104] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1486__I0 (.I(\mod.buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__A1 (.I(\mod.buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__I1 (.I(\mod.buffer[134] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__I0 (.I(\mod.buffer[134] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1421__A1 (.I(\mod.buffer[134] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__I1 (.I(\mod.buffer[136] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__I0 (.I(\mod.buffer[136] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A1 (.I(\mod.buffer[136] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__I1 (.I(\mod.buffer[139] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A1 (.I(\mod.buffer[139] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__A1 (.I(\mod.buffer[139] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__I (.I(\mod.buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0908__I (.I(\mod.buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__I0 (.I(\mod.buffer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__I1 (.I(\mod.buffer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__I0 (.I(\mod.buffer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__I1 (.I(\mod.buffer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__I0 (.I(\mod.buffer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__I1 (.I(\mod.buffer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__I (.I(\mod.buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0982__I (.I(\mod.buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0945__I (.I(\mod.buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__I (.I(\mod.buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__I0 (.I(\mod.buffer[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__I1 (.I(\mod.buffer[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__I0 (.I(\mod.buffer[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__I1 (.I(\mod.buffer[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1049__I (.I(\mod.buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1033__I (.I(\mod.buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1011__I (.I(\mod.buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0964__I (.I(\mod.buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__I0 (.I(\mod.buffer[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__I1 (.I(\mod.buffer[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__I0 (.I(\mod.buffer[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__I1 (.I(\mod.buffer[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__I0 (.I(\mod.buffer[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__I1 (.I(\mod.buffer[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1147__I (.I(\mod.buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__I (.I(\mod.buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__I (.I(\mod.buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__I (.I(\mod.buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I0 (.I(\mod.buffer[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__I1 (.I(\mod.buffer[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0904__I (.I(\mod.buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0885__A2 (.I(\mod.buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__I0 (.I(\mod.buffer[96] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__I1 (.I(\mod.buffer[96] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0917__I (.I(\mod.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0888__A2 (.I(\mod.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0881__I (.I(\mod.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__I (.I(\mod.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0887__I (.I(\mod.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0946__A3 (.I(\mod.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0914__I (.I(\mod.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0900__I (.I(\mod.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0892__I (.I(\mod.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0885__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__B2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1048__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__CLK (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__CLK (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout15_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout16_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__CLK (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__CLK (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__CLK (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__CLK (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__CLK (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__CLK (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__CLK (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__CLK (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__CLK (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__CLK (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout19_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout17_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__CLK (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__CLK (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__CLK (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__CLK (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__CLK (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout24_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__CLK (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout23_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout26_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__CLK (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__CLK (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__CLK (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout27_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__CLK (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__CLK (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__CLK (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__CLK (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__CLK (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__CLK (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1758 ();
 assign io_oeb[0] = net75;
 assign io_oeb[10] = net85;
 assign io_oeb[11] = net86;
 assign io_oeb[12] = net87;
 assign io_oeb[13] = net88;
 assign io_oeb[14] = net89;
 assign io_oeb[15] = net90;
 assign io_oeb[16] = net91;
 assign io_oeb[17] = net92;
 assign io_oeb[18] = net93;
 assign io_oeb[19] = net94;
 assign io_oeb[1] = net76;
 assign io_oeb[20] = net95;
 assign io_oeb[21] = net96;
 assign io_oeb[22] = net97;
 assign io_oeb[23] = net98;
 assign io_oeb[24] = net99;
 assign io_oeb[25] = net100;
 assign io_oeb[26] = net101;
 assign io_oeb[27] = net102;
 assign io_oeb[28] = net103;
 assign io_oeb[29] = net104;
 assign io_oeb[2] = net77;
 assign io_oeb[30] = net105;
 assign io_oeb[31] = net106;
 assign io_oeb[32] = net107;
 assign io_oeb[33] = net108;
 assign io_oeb[34] = net109;
 assign io_oeb[35] = net110;
 assign io_oeb[36] = net111;
 assign io_oeb[37] = net112;
 assign io_oeb[3] = net78;
 assign io_oeb[4] = net79;
 assign io_oeb[5] = net80;
 assign io_oeb[6] = net81;
 assign io_oeb[7] = net82;
 assign io_oeb[8] = net83;
 assign io_oeb[9] = net84;
 assign io_out[0] = net113;
 assign io_out[10] = net123;
 assign io_out[11] = net124;
 assign io_out[12] = net125;
 assign io_out[13] = net126;
 assign io_out[14] = net127;
 assign io_out[15] = net128;
 assign io_out[1] = net114;
 assign io_out[24] = net129;
 assign io_out[25] = net130;
 assign io_out[26] = net131;
 assign io_out[27] = net132;
 assign io_out[28] = net133;
 assign io_out[29] = net134;
 assign io_out[2] = net115;
 assign io_out[30] = net135;
 assign io_out[31] = net136;
 assign io_out[32] = net137;
 assign io_out[33] = net138;
 assign io_out[34] = net139;
 assign io_out[35] = net140;
 assign io_out[36] = net141;
 assign io_out[37] = net142;
 assign io_out[3] = net116;
 assign io_out[4] = net117;
 assign io_out[5] = net118;
 assign io_out[6] = net119;
 assign io_out[7] = net120;
 assign io_out[8] = net121;
 assign io_out[9] = net122;
 assign la_data_out[0] = net143;
 assign la_data_out[10] = net153;
 assign la_data_out[11] = net154;
 assign la_data_out[12] = net155;
 assign la_data_out[13] = net156;
 assign la_data_out[14] = net157;
 assign la_data_out[15] = net158;
 assign la_data_out[16] = net159;
 assign la_data_out[17] = net160;
 assign la_data_out[18] = net161;
 assign la_data_out[19] = net162;
 assign la_data_out[1] = net144;
 assign la_data_out[20] = net163;
 assign la_data_out[21] = net164;
 assign la_data_out[22] = net165;
 assign la_data_out[23] = net166;
 assign la_data_out[24] = net167;
 assign la_data_out[25] = net168;
 assign la_data_out[26] = net169;
 assign la_data_out[27] = net170;
 assign la_data_out[28] = net171;
 assign la_data_out[29] = net172;
 assign la_data_out[2] = net145;
 assign la_data_out[30] = net173;
 assign la_data_out[31] = net174;
 assign la_data_out[32] = net175;
 assign la_data_out[33] = net176;
 assign la_data_out[34] = net177;
 assign la_data_out[35] = net178;
 assign la_data_out[36] = net179;
 assign la_data_out[37] = net180;
 assign la_data_out[38] = net181;
 assign la_data_out[39] = net182;
 assign la_data_out[3] = net146;
 assign la_data_out[40] = net183;
 assign la_data_out[41] = net184;
 assign la_data_out[42] = net185;
 assign la_data_out[43] = net186;
 assign la_data_out[44] = net187;
 assign la_data_out[45] = net188;
 assign la_data_out[46] = net189;
 assign la_data_out[47] = net190;
 assign la_data_out[48] = net191;
 assign la_data_out[49] = net192;
 assign la_data_out[4] = net147;
 assign la_data_out[50] = net193;
 assign la_data_out[51] = net194;
 assign la_data_out[52] = net195;
 assign la_data_out[53] = net196;
 assign la_data_out[54] = net197;
 assign la_data_out[55] = net198;
 assign la_data_out[56] = net199;
 assign la_data_out[57] = net200;
 assign la_data_out[58] = net201;
 assign la_data_out[59] = net202;
 assign la_data_out[5] = net148;
 assign la_data_out[60] = net203;
 assign la_data_out[61] = net204;
 assign la_data_out[62] = net205;
 assign la_data_out[63] = net206;
 assign la_data_out[6] = net149;
 assign la_data_out[7] = net150;
 assign la_data_out[8] = net151;
 assign la_data_out[9] = net152;
 assign user_irq[0] = net207;
 assign user_irq[1] = net208;
 assign user_irq[2] = net209;
 assign wbs_ack_o = net210;
 assign wbs_dat_o[0] = net211;
 assign wbs_dat_o[10] = net221;
 assign wbs_dat_o[11] = net222;
 assign wbs_dat_o[12] = net223;
 assign wbs_dat_o[13] = net224;
 assign wbs_dat_o[14] = net225;
 assign wbs_dat_o[15] = net226;
 assign wbs_dat_o[16] = net227;
 assign wbs_dat_o[17] = net228;
 assign wbs_dat_o[18] = net229;
 assign wbs_dat_o[19] = net230;
 assign wbs_dat_o[1] = net212;
 assign wbs_dat_o[20] = net231;
 assign wbs_dat_o[21] = net232;
 assign wbs_dat_o[22] = net233;
 assign wbs_dat_o[23] = net234;
 assign wbs_dat_o[24] = net235;
 assign wbs_dat_o[25] = net236;
 assign wbs_dat_o[26] = net237;
 assign wbs_dat_o[27] = net238;
 assign wbs_dat_o[28] = net239;
 assign wbs_dat_o[29] = net240;
 assign wbs_dat_o[2] = net213;
 assign wbs_dat_o[30] = net241;
 assign wbs_dat_o[31] = net242;
 assign wbs_dat_o[3] = net214;
 assign wbs_dat_o[4] = net215;
 assign wbs_dat_o[5] = net216;
 assign wbs_dat_o[6] = net217;
 assign wbs_dat_o[7] = net218;
 assign wbs_dat_o[8] = net219;
 assign wbs_dat_o[9] = net220;
endmodule

