magic
tech gf180mcuC
magscale 1 5
timestamp 1670248760
<< obsm1 >>
rect 672 911 99288 98422
<< metal2 >>
rect 672 99600 728 99900
rect 1680 99600 1736 99900
rect 2688 99600 2744 99900
rect 3696 99600 3752 99900
rect 4704 99600 4760 99900
rect 5712 99600 5768 99900
rect 6720 99600 6776 99900
rect 7392 99600 7448 99900
rect 8400 99600 8456 99900
rect 9408 99600 9464 99900
rect 10416 99600 10472 99900
rect 11424 99600 11480 99900
rect 12432 99600 12488 99900
rect 13440 99600 13496 99900
rect 14112 99600 14168 99900
rect 15120 99600 15176 99900
rect 16128 99600 16184 99900
rect 17136 99600 17192 99900
rect 18144 99600 18200 99900
rect 19152 99600 19208 99900
rect 20160 99600 20216 99900
rect 21168 99600 21224 99900
rect 21840 99600 21896 99900
rect 22848 99600 22904 99900
rect 23856 99600 23912 99900
rect 24864 99600 24920 99900
rect 25872 99600 25928 99900
rect 26880 99600 26936 99900
rect 27888 99600 27944 99900
rect 28560 99600 28616 99900
rect 29568 99600 29624 99900
rect 30576 99600 30632 99900
rect 31584 99600 31640 99900
rect 32592 99600 32648 99900
rect 33600 99600 33656 99900
rect 34608 99600 34664 99900
rect 35616 99600 35672 99900
rect 36288 99600 36344 99900
rect 37296 99600 37352 99900
rect 38304 99600 38360 99900
rect 39312 99600 39368 99900
rect 40320 99600 40376 99900
rect 41328 99600 41384 99900
rect 42336 99600 42392 99900
rect 43008 99600 43064 99900
rect 44016 99600 44072 99900
rect 45024 99600 45080 99900
rect 46032 99600 46088 99900
rect 47040 99600 47096 99900
rect 48048 99600 48104 99900
rect 49056 99600 49112 99900
rect 49728 99600 49784 99900
rect 50736 99600 50792 99900
rect 51744 99600 51800 99900
rect 52752 99600 52808 99900
rect 53760 99600 53816 99900
rect 54768 99600 54824 99900
rect 55776 99600 55832 99900
rect 56784 99600 56840 99900
rect 57456 99600 57512 99900
rect 58464 99600 58520 99900
rect 59472 99600 59528 99900
rect 60480 99600 60536 99900
rect 61488 99600 61544 99900
rect 62496 99600 62552 99900
rect 63504 99600 63560 99900
rect 64176 99600 64232 99900
rect 65184 99600 65240 99900
rect 66192 99600 66248 99900
rect 67200 99600 67256 99900
rect 68208 99600 68264 99900
rect 69216 99600 69272 99900
rect 70224 99600 70280 99900
rect 71232 99600 71288 99900
rect 71904 99600 71960 99900
rect 72912 99600 72968 99900
rect 73920 99600 73976 99900
rect 74928 99600 74984 99900
rect 75936 99600 75992 99900
rect 76944 99600 77000 99900
rect 77952 99600 78008 99900
rect 78624 99600 78680 99900
rect 79632 99600 79688 99900
rect 80640 99600 80696 99900
rect 81648 99600 81704 99900
rect 82656 99600 82712 99900
rect 83664 99600 83720 99900
rect 84672 99600 84728 99900
rect 85680 99600 85736 99900
rect 86352 99600 86408 99900
rect 87360 99600 87416 99900
rect 88368 99600 88424 99900
rect 89376 99600 89432 99900
rect 90384 99600 90440 99900
rect 91392 99600 91448 99900
rect 92400 99600 92456 99900
rect 93072 99600 93128 99900
rect 94080 99600 94136 99900
rect 95088 99600 95144 99900
rect 96096 99600 96152 99900
rect 97104 99600 97160 99900
rect 98112 99600 98168 99900
rect 99120 99600 99176 99900
rect 99792 99600 99848 99900
rect 0 100 56 400
rect 672 100 728 400
rect 1680 100 1736 400
rect 2688 100 2744 400
rect 3696 100 3752 400
rect 4704 100 4760 400
rect 5712 100 5768 400
rect 6720 100 6776 400
rect 7392 100 7448 400
rect 8400 100 8456 400
rect 9408 100 9464 400
rect 10416 100 10472 400
rect 11424 100 11480 400
rect 12432 100 12488 400
rect 13440 100 13496 400
rect 14112 100 14168 400
rect 15120 100 15176 400
rect 16128 100 16184 400
rect 17136 100 17192 400
rect 18144 100 18200 400
rect 19152 100 19208 400
rect 20160 100 20216 400
rect 21168 100 21224 400
rect 21840 100 21896 400
rect 22848 100 22904 400
rect 23856 100 23912 400
rect 24864 100 24920 400
rect 25872 100 25928 400
rect 26880 100 26936 400
rect 27888 100 27944 400
rect 28560 100 28616 400
rect 29568 100 29624 400
rect 30576 100 30632 400
rect 31584 100 31640 400
rect 32592 100 32648 400
rect 33600 100 33656 400
rect 34608 100 34664 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 37296 100 37352 400
rect 38304 100 38360 400
rect 39312 100 39368 400
rect 40320 100 40376 400
rect 41328 100 41384 400
rect 42336 100 42392 400
rect 43008 100 43064 400
rect 44016 100 44072 400
rect 45024 100 45080 400
rect 46032 100 46088 400
rect 47040 100 47096 400
rect 48048 100 48104 400
rect 49056 100 49112 400
rect 50064 100 50120 400
rect 50736 100 50792 400
rect 51744 100 51800 400
rect 52752 100 52808 400
rect 53760 100 53816 400
rect 54768 100 54824 400
rect 55776 100 55832 400
rect 56784 100 56840 400
rect 57456 100 57512 400
rect 58464 100 58520 400
rect 59472 100 59528 400
rect 60480 100 60536 400
rect 61488 100 61544 400
rect 62496 100 62552 400
rect 63504 100 63560 400
rect 64176 100 64232 400
rect 65184 100 65240 400
rect 66192 100 66248 400
rect 67200 100 67256 400
rect 68208 100 68264 400
rect 69216 100 69272 400
rect 70224 100 70280 400
rect 71232 100 71288 400
rect 71904 100 71960 400
rect 72912 100 72968 400
rect 73920 100 73976 400
rect 74928 100 74984 400
rect 75936 100 75992 400
rect 76944 100 77000 400
rect 77952 100 78008 400
rect 78624 100 78680 400
rect 79632 100 79688 400
rect 80640 100 80696 400
rect 81648 100 81704 400
rect 82656 100 82712 400
rect 83664 100 83720 400
rect 84672 100 84728 400
rect 85680 100 85736 400
rect 86352 100 86408 400
rect 87360 100 87416 400
rect 88368 100 88424 400
rect 89376 100 89432 400
rect 90384 100 90440 400
rect 91392 100 91448 400
rect 92400 100 92456 400
rect 93072 100 93128 400
rect 94080 100 94136 400
rect 95088 100 95144 400
rect 96096 100 96152 400
rect 97104 100 97160 400
rect 98112 100 98168 400
rect 99120 100 99176 400
<< obsm2 >>
rect 14 99570 642 99839
rect 758 99570 1650 99839
rect 1766 99570 2658 99839
rect 2774 99570 3666 99839
rect 3782 99570 4674 99839
rect 4790 99570 5682 99839
rect 5798 99570 6690 99839
rect 6806 99570 7362 99839
rect 7478 99570 8370 99839
rect 8486 99570 9378 99839
rect 9494 99570 10386 99839
rect 10502 99570 11394 99839
rect 11510 99570 12402 99839
rect 12518 99570 13410 99839
rect 13526 99570 14082 99839
rect 14198 99570 15090 99839
rect 15206 99570 16098 99839
rect 16214 99570 17106 99839
rect 17222 99570 18114 99839
rect 18230 99570 19122 99839
rect 19238 99570 20130 99839
rect 20246 99570 21138 99839
rect 21254 99570 21810 99839
rect 21926 99570 22818 99839
rect 22934 99570 23826 99839
rect 23942 99570 24834 99839
rect 24950 99570 25842 99839
rect 25958 99570 26850 99839
rect 26966 99570 27858 99839
rect 27974 99570 28530 99839
rect 28646 99570 29538 99839
rect 29654 99570 30546 99839
rect 30662 99570 31554 99839
rect 31670 99570 32562 99839
rect 32678 99570 33570 99839
rect 33686 99570 34578 99839
rect 34694 99570 35586 99839
rect 35702 99570 36258 99839
rect 36374 99570 37266 99839
rect 37382 99570 38274 99839
rect 38390 99570 39282 99839
rect 39398 99570 40290 99839
rect 40406 99570 41298 99839
rect 41414 99570 42306 99839
rect 42422 99570 42978 99839
rect 43094 99570 43986 99839
rect 44102 99570 44994 99839
rect 45110 99570 46002 99839
rect 46118 99570 47010 99839
rect 47126 99570 48018 99839
rect 48134 99570 49026 99839
rect 49142 99570 49698 99839
rect 49814 99570 50706 99839
rect 50822 99570 51714 99839
rect 51830 99570 52722 99839
rect 52838 99570 53730 99839
rect 53846 99570 54738 99839
rect 54854 99570 55746 99839
rect 55862 99570 56754 99839
rect 56870 99570 57426 99839
rect 57542 99570 58434 99839
rect 58550 99570 59442 99839
rect 59558 99570 60450 99839
rect 60566 99570 61458 99839
rect 61574 99570 62466 99839
rect 62582 99570 63474 99839
rect 63590 99570 64146 99839
rect 64262 99570 65154 99839
rect 65270 99570 66162 99839
rect 66278 99570 67170 99839
rect 67286 99570 68178 99839
rect 68294 99570 69186 99839
rect 69302 99570 70194 99839
rect 70310 99570 71202 99839
rect 71318 99570 71874 99839
rect 71990 99570 72882 99839
rect 72998 99570 73890 99839
rect 74006 99570 74898 99839
rect 75014 99570 75906 99839
rect 76022 99570 76914 99839
rect 77030 99570 77922 99839
rect 78038 99570 78594 99839
rect 78710 99570 79602 99839
rect 79718 99570 80610 99839
rect 80726 99570 81618 99839
rect 81734 99570 82626 99839
rect 82742 99570 83634 99839
rect 83750 99570 84642 99839
rect 84758 99570 85650 99839
rect 85766 99570 86322 99839
rect 86438 99570 87330 99839
rect 87446 99570 88338 99839
rect 88454 99570 89346 99839
rect 89462 99570 90354 99839
rect 90470 99570 91362 99839
rect 91478 99570 92370 99839
rect 92486 99570 93042 99839
rect 93158 99570 94050 99839
rect 94166 99570 95058 99839
rect 95174 99570 96066 99839
rect 96182 99570 97074 99839
rect 97190 99570 98082 99839
rect 98198 99570 99090 99839
rect 14 430 99162 99570
rect 86 400 642 430
rect 758 400 1650 430
rect 1766 400 2658 430
rect 2774 400 3666 430
rect 3782 400 4674 430
rect 4790 400 5682 430
rect 5798 400 6690 430
rect 6806 400 7362 430
rect 7478 400 8370 430
rect 8486 400 9378 430
rect 9494 400 10386 430
rect 10502 400 11394 430
rect 11510 400 12402 430
rect 12518 400 13410 430
rect 13526 400 14082 430
rect 14198 400 15090 430
rect 15206 400 16098 430
rect 16214 400 17106 430
rect 17222 400 18114 430
rect 18230 400 19122 430
rect 19238 400 20130 430
rect 20246 400 21138 430
rect 21254 400 21810 430
rect 21926 400 22818 430
rect 22934 400 23826 430
rect 23942 400 24834 430
rect 24950 400 25842 430
rect 25958 400 26850 430
rect 26966 400 27858 430
rect 27974 400 28530 430
rect 28646 400 29538 430
rect 29654 400 30546 430
rect 30662 400 31554 430
rect 31670 400 32562 430
rect 32678 400 33570 430
rect 33686 400 34578 430
rect 34694 400 35586 430
rect 35702 400 36258 430
rect 36374 400 37266 430
rect 37382 400 38274 430
rect 38390 400 39282 430
rect 39398 400 40290 430
rect 40406 400 41298 430
rect 41414 400 42306 430
rect 42422 400 42978 430
rect 43094 400 43986 430
rect 44102 400 44994 430
rect 45110 400 46002 430
rect 46118 400 47010 430
rect 47126 400 48018 430
rect 48134 400 49026 430
rect 49142 400 50034 430
rect 50150 400 50706 430
rect 50822 400 51714 430
rect 51830 400 52722 430
rect 52838 400 53730 430
rect 53846 400 54738 430
rect 54854 400 55746 430
rect 55862 400 56754 430
rect 56870 400 57426 430
rect 57542 400 58434 430
rect 58550 400 59442 430
rect 59558 400 60450 430
rect 60566 400 61458 430
rect 61574 400 62466 430
rect 62582 400 63474 430
rect 63590 400 64146 430
rect 64262 400 65154 430
rect 65270 400 66162 430
rect 66278 400 67170 430
rect 67286 400 68178 430
rect 68294 400 69186 430
rect 69302 400 70194 430
rect 70310 400 71202 430
rect 71318 400 71874 430
rect 71990 400 72882 430
rect 72998 400 73890 430
rect 74006 400 74898 430
rect 75014 400 75906 430
rect 76022 400 76914 430
rect 77030 400 77922 430
rect 78038 400 78594 430
rect 78710 400 79602 430
rect 79718 400 80610 430
rect 80726 400 81618 430
rect 81734 400 82626 430
rect 82742 400 83634 430
rect 83750 400 84642 430
rect 84758 400 85650 430
rect 85766 400 86322 430
rect 86438 400 87330 430
rect 87446 400 88338 430
rect 88454 400 89346 430
rect 89462 400 90354 430
rect 90470 400 91362 430
rect 91478 400 92370 430
rect 92486 400 93042 430
rect 93158 400 94050 430
rect 94166 400 95058 430
rect 95174 400 96066 430
rect 96182 400 97074 430
rect 97190 400 98082 430
rect 98198 400 99090 430
<< metal3 >>
rect 100 99792 400 99848
rect 100 99120 400 99176
rect 99600 99120 99900 99176
rect 100 98112 400 98168
rect 99600 98112 99900 98168
rect 100 97104 400 97160
rect 99600 97104 99900 97160
rect 100 96096 400 96152
rect 99600 96096 99900 96152
rect 100 95088 400 95144
rect 99600 95088 99900 95144
rect 100 94080 400 94136
rect 99600 94080 99900 94136
rect 100 93072 400 93128
rect 99600 93072 99900 93128
rect 100 92400 400 92456
rect 99600 92400 99900 92456
rect 100 91392 400 91448
rect 99600 91392 99900 91448
rect 100 90384 400 90440
rect 99600 90384 99900 90440
rect 100 89376 400 89432
rect 99600 89376 99900 89432
rect 100 88368 400 88424
rect 99600 88368 99900 88424
rect 100 87360 400 87416
rect 99600 87360 99900 87416
rect 100 86352 400 86408
rect 99600 86352 99900 86408
rect 100 85680 400 85736
rect 99600 85680 99900 85736
rect 100 84672 400 84728
rect 99600 84672 99900 84728
rect 100 83664 400 83720
rect 99600 83664 99900 83720
rect 100 82656 400 82712
rect 99600 82656 99900 82712
rect 100 81648 400 81704
rect 99600 81648 99900 81704
rect 100 80640 400 80696
rect 99600 80640 99900 80696
rect 100 79632 400 79688
rect 99600 79632 99900 79688
rect 100 78624 400 78680
rect 99600 78624 99900 78680
rect 100 77952 400 78008
rect 99600 77952 99900 78008
rect 100 76944 400 77000
rect 99600 76944 99900 77000
rect 100 75936 400 75992
rect 99600 75936 99900 75992
rect 100 74928 400 74984
rect 99600 74928 99900 74984
rect 100 73920 400 73976
rect 99600 73920 99900 73976
rect 100 72912 400 72968
rect 99600 72912 99900 72968
rect 100 71904 400 71960
rect 99600 71904 99900 71960
rect 100 71232 400 71288
rect 99600 71232 99900 71288
rect 100 70224 400 70280
rect 99600 70224 99900 70280
rect 100 69216 400 69272
rect 99600 69216 99900 69272
rect 100 68208 400 68264
rect 99600 68208 99900 68264
rect 100 67200 400 67256
rect 99600 67200 99900 67256
rect 100 66192 400 66248
rect 99600 66192 99900 66248
rect 100 65184 400 65240
rect 99600 65184 99900 65240
rect 100 64176 400 64232
rect 99600 64176 99900 64232
rect 100 63504 400 63560
rect 99600 63504 99900 63560
rect 100 62496 400 62552
rect 99600 62496 99900 62552
rect 100 61488 400 61544
rect 99600 61488 99900 61544
rect 100 60480 400 60536
rect 99600 60480 99900 60536
rect 100 59472 400 59528
rect 99600 59472 99900 59528
rect 100 58464 400 58520
rect 99600 58464 99900 58520
rect 100 57456 400 57512
rect 99600 57456 99900 57512
rect 100 56784 400 56840
rect 99600 56784 99900 56840
rect 100 55776 400 55832
rect 99600 55776 99900 55832
rect 100 54768 400 54824
rect 99600 54768 99900 54824
rect 100 53760 400 53816
rect 99600 53760 99900 53816
rect 100 52752 400 52808
rect 99600 52752 99900 52808
rect 100 51744 400 51800
rect 99600 51744 99900 51800
rect 100 50736 400 50792
rect 99600 50736 99900 50792
rect 99600 50064 99900 50120
rect 100 49728 400 49784
rect 100 49056 400 49112
rect 99600 49056 99900 49112
rect 100 48048 400 48104
rect 99600 48048 99900 48104
rect 100 47040 400 47096
rect 99600 47040 99900 47096
rect 100 46032 400 46088
rect 99600 46032 99900 46088
rect 100 45024 400 45080
rect 99600 45024 99900 45080
rect 100 44016 400 44072
rect 99600 44016 99900 44072
rect 100 43008 400 43064
rect 99600 43008 99900 43064
rect 100 42336 400 42392
rect 99600 42336 99900 42392
rect 100 41328 400 41384
rect 99600 41328 99900 41384
rect 100 40320 400 40376
rect 99600 40320 99900 40376
rect 100 39312 400 39368
rect 99600 39312 99900 39368
rect 100 38304 400 38360
rect 99600 38304 99900 38360
rect 100 37296 400 37352
rect 99600 37296 99900 37352
rect 100 36288 400 36344
rect 99600 36288 99900 36344
rect 100 35616 400 35672
rect 99600 35616 99900 35672
rect 100 34608 400 34664
rect 99600 34608 99900 34664
rect 100 33600 400 33656
rect 99600 33600 99900 33656
rect 100 32592 400 32648
rect 99600 32592 99900 32648
rect 100 31584 400 31640
rect 99600 31584 99900 31640
rect 100 30576 400 30632
rect 99600 30576 99900 30632
rect 100 29568 400 29624
rect 99600 29568 99900 29624
rect 100 28560 400 28616
rect 99600 28560 99900 28616
rect 100 27888 400 27944
rect 99600 27888 99900 27944
rect 100 26880 400 26936
rect 99600 26880 99900 26936
rect 100 25872 400 25928
rect 99600 25872 99900 25928
rect 100 24864 400 24920
rect 99600 24864 99900 24920
rect 100 23856 400 23912
rect 99600 23856 99900 23912
rect 100 22848 400 22904
rect 99600 22848 99900 22904
rect 100 21840 400 21896
rect 99600 21840 99900 21896
rect 100 21168 400 21224
rect 99600 21168 99900 21224
rect 100 20160 400 20216
rect 99600 20160 99900 20216
rect 100 19152 400 19208
rect 99600 19152 99900 19208
rect 100 18144 400 18200
rect 99600 18144 99900 18200
rect 100 17136 400 17192
rect 99600 17136 99900 17192
rect 100 16128 400 16184
rect 99600 16128 99900 16184
rect 100 15120 400 15176
rect 99600 15120 99900 15176
rect 100 14112 400 14168
rect 99600 14112 99900 14168
rect 100 13440 400 13496
rect 99600 13440 99900 13496
rect 100 12432 400 12488
rect 99600 12432 99900 12488
rect 100 11424 400 11480
rect 99600 11424 99900 11480
rect 100 10416 400 10472
rect 99600 10416 99900 10472
rect 100 9408 400 9464
rect 99600 9408 99900 9464
rect 100 8400 400 8456
rect 99600 8400 99900 8456
rect 100 7392 400 7448
rect 99600 7392 99900 7448
rect 100 6720 400 6776
rect 99600 6720 99900 6776
rect 100 5712 400 5768
rect 99600 5712 99900 5768
rect 100 4704 400 4760
rect 99600 4704 99900 4760
rect 100 3696 400 3752
rect 99600 3696 99900 3752
rect 100 2688 400 2744
rect 99600 2688 99900 2744
rect 100 1680 400 1736
rect 99600 1680 99900 1736
rect 100 672 400 728
rect 99600 672 99900 728
rect 99600 0 99900 56
<< obsm3 >>
rect 9 99762 70 99834
rect 430 99762 99600 99834
rect 9 99206 99600 99762
rect 9 99090 70 99206
rect 430 99090 99570 99206
rect 9 98198 99600 99090
rect 9 98082 70 98198
rect 430 98082 99570 98198
rect 9 97190 99600 98082
rect 9 97074 70 97190
rect 430 97074 99570 97190
rect 9 96182 99600 97074
rect 9 96066 70 96182
rect 430 96066 99570 96182
rect 9 95174 99600 96066
rect 9 95058 70 95174
rect 430 95058 99570 95174
rect 9 94166 99600 95058
rect 9 94050 70 94166
rect 430 94050 99570 94166
rect 9 93158 99600 94050
rect 9 93042 70 93158
rect 430 93042 99570 93158
rect 9 92486 99600 93042
rect 9 92370 70 92486
rect 430 92370 99570 92486
rect 9 91478 99600 92370
rect 9 91362 70 91478
rect 430 91362 99570 91478
rect 9 90470 99600 91362
rect 9 90354 70 90470
rect 430 90354 99570 90470
rect 9 89462 99600 90354
rect 9 89346 70 89462
rect 430 89346 99570 89462
rect 9 88454 99600 89346
rect 9 88338 70 88454
rect 430 88338 99570 88454
rect 9 87446 99600 88338
rect 9 87330 70 87446
rect 430 87330 99570 87446
rect 9 86438 99600 87330
rect 9 86322 70 86438
rect 430 86322 99570 86438
rect 9 85766 99600 86322
rect 9 85650 70 85766
rect 430 85650 99570 85766
rect 9 84758 99600 85650
rect 9 84642 70 84758
rect 430 84642 99570 84758
rect 9 83750 99600 84642
rect 9 83634 70 83750
rect 430 83634 99570 83750
rect 9 82742 99600 83634
rect 9 82626 70 82742
rect 430 82626 99570 82742
rect 9 81734 99600 82626
rect 9 81618 70 81734
rect 430 81618 99570 81734
rect 9 80726 99600 81618
rect 9 80610 70 80726
rect 430 80610 99570 80726
rect 9 79718 99600 80610
rect 9 79602 70 79718
rect 430 79602 99570 79718
rect 9 78710 99600 79602
rect 9 78594 70 78710
rect 430 78594 99570 78710
rect 9 78038 99600 78594
rect 9 77922 70 78038
rect 430 77922 99570 78038
rect 9 77030 99600 77922
rect 9 76914 70 77030
rect 430 76914 99570 77030
rect 9 76022 99600 76914
rect 9 75906 70 76022
rect 430 75906 99570 76022
rect 9 75014 99600 75906
rect 9 74898 70 75014
rect 430 74898 99570 75014
rect 9 74006 99600 74898
rect 9 73890 70 74006
rect 430 73890 99570 74006
rect 9 72998 99600 73890
rect 9 72882 70 72998
rect 430 72882 99570 72998
rect 9 71990 99600 72882
rect 9 71874 70 71990
rect 430 71874 99570 71990
rect 9 71318 99600 71874
rect 9 71202 70 71318
rect 430 71202 99570 71318
rect 9 70310 99600 71202
rect 9 70194 70 70310
rect 430 70194 99570 70310
rect 9 69302 99600 70194
rect 9 69186 70 69302
rect 430 69186 99570 69302
rect 9 68294 99600 69186
rect 9 68178 70 68294
rect 430 68178 99570 68294
rect 9 67286 99600 68178
rect 9 67170 70 67286
rect 430 67170 99570 67286
rect 9 66278 99600 67170
rect 9 66162 70 66278
rect 430 66162 99570 66278
rect 9 65270 99600 66162
rect 9 65154 70 65270
rect 430 65154 99570 65270
rect 9 64262 99600 65154
rect 9 64146 70 64262
rect 430 64146 99570 64262
rect 9 63590 99600 64146
rect 9 63474 70 63590
rect 430 63474 99570 63590
rect 9 62582 99600 63474
rect 9 62466 70 62582
rect 430 62466 99570 62582
rect 9 61574 99600 62466
rect 9 61458 70 61574
rect 430 61458 99570 61574
rect 9 60566 99600 61458
rect 9 60450 70 60566
rect 430 60450 99570 60566
rect 9 59558 99600 60450
rect 9 59442 70 59558
rect 430 59442 99570 59558
rect 9 58550 99600 59442
rect 9 58434 70 58550
rect 430 58434 99570 58550
rect 9 57542 99600 58434
rect 9 57426 70 57542
rect 430 57426 99570 57542
rect 9 56870 99600 57426
rect 9 56754 70 56870
rect 430 56754 99570 56870
rect 9 55862 99600 56754
rect 9 55746 70 55862
rect 430 55746 99570 55862
rect 9 54854 99600 55746
rect 9 54738 70 54854
rect 430 54738 99570 54854
rect 9 53846 99600 54738
rect 9 53730 70 53846
rect 430 53730 99570 53846
rect 9 52838 99600 53730
rect 9 52722 70 52838
rect 430 52722 99570 52838
rect 9 51830 99600 52722
rect 9 51714 70 51830
rect 430 51714 99570 51830
rect 9 50822 99600 51714
rect 9 50706 70 50822
rect 430 50706 99570 50822
rect 9 50150 99600 50706
rect 9 50034 99570 50150
rect 9 49814 99600 50034
rect 9 49698 70 49814
rect 430 49698 99600 49814
rect 9 49142 99600 49698
rect 9 49026 70 49142
rect 430 49026 99570 49142
rect 9 48134 99600 49026
rect 9 48018 70 48134
rect 430 48018 99570 48134
rect 9 47126 99600 48018
rect 9 47010 70 47126
rect 430 47010 99570 47126
rect 9 46118 99600 47010
rect 9 46002 70 46118
rect 430 46002 99570 46118
rect 9 45110 99600 46002
rect 9 44994 70 45110
rect 430 44994 99570 45110
rect 9 44102 99600 44994
rect 9 43986 70 44102
rect 430 43986 99570 44102
rect 9 43094 99600 43986
rect 9 42978 70 43094
rect 430 42978 99570 43094
rect 9 42422 99600 42978
rect 9 42306 70 42422
rect 430 42306 99570 42422
rect 9 41414 99600 42306
rect 9 41298 70 41414
rect 430 41298 99570 41414
rect 9 40406 99600 41298
rect 9 40290 70 40406
rect 430 40290 99570 40406
rect 9 39398 99600 40290
rect 9 39282 70 39398
rect 430 39282 99570 39398
rect 9 38390 99600 39282
rect 9 38274 70 38390
rect 430 38274 99570 38390
rect 9 37382 99600 38274
rect 9 37266 70 37382
rect 430 37266 99570 37382
rect 9 36374 99600 37266
rect 9 36258 70 36374
rect 430 36258 99570 36374
rect 9 35702 99600 36258
rect 9 35586 70 35702
rect 430 35586 99570 35702
rect 9 34694 99600 35586
rect 9 34578 70 34694
rect 430 34578 99570 34694
rect 9 33686 99600 34578
rect 9 33570 70 33686
rect 430 33570 99570 33686
rect 9 32678 99600 33570
rect 9 32562 70 32678
rect 430 32562 99570 32678
rect 9 31670 99600 32562
rect 9 31554 70 31670
rect 430 31554 99570 31670
rect 9 30662 99600 31554
rect 9 30546 70 30662
rect 430 30546 99570 30662
rect 9 29654 99600 30546
rect 9 29538 70 29654
rect 430 29538 99570 29654
rect 9 28646 99600 29538
rect 9 28530 70 28646
rect 430 28530 99570 28646
rect 9 27974 99600 28530
rect 9 27858 70 27974
rect 430 27858 99570 27974
rect 9 26966 99600 27858
rect 9 26850 70 26966
rect 430 26850 99570 26966
rect 9 25958 99600 26850
rect 9 25842 70 25958
rect 430 25842 99570 25958
rect 9 24950 99600 25842
rect 9 24834 70 24950
rect 430 24834 99570 24950
rect 9 23942 99600 24834
rect 9 23826 70 23942
rect 430 23826 99570 23942
rect 9 22934 99600 23826
rect 9 22818 70 22934
rect 430 22818 99570 22934
rect 9 21926 99600 22818
rect 9 21810 70 21926
rect 430 21810 99570 21926
rect 9 21254 99600 21810
rect 9 21138 70 21254
rect 430 21138 99570 21254
rect 9 20246 99600 21138
rect 9 20130 70 20246
rect 430 20130 99570 20246
rect 9 19238 99600 20130
rect 9 19122 70 19238
rect 430 19122 99570 19238
rect 9 18230 99600 19122
rect 9 18114 70 18230
rect 430 18114 99570 18230
rect 9 17222 99600 18114
rect 9 17106 70 17222
rect 430 17106 99570 17222
rect 9 16214 99600 17106
rect 9 16098 70 16214
rect 430 16098 99570 16214
rect 9 15206 99600 16098
rect 9 15090 70 15206
rect 430 15090 99570 15206
rect 9 14198 99600 15090
rect 9 14082 70 14198
rect 430 14082 99570 14198
rect 9 13526 99600 14082
rect 9 13410 70 13526
rect 430 13410 99570 13526
rect 9 12518 99600 13410
rect 9 12402 70 12518
rect 430 12402 99570 12518
rect 9 11510 99600 12402
rect 9 11394 70 11510
rect 430 11394 99570 11510
rect 9 10502 99600 11394
rect 9 10386 70 10502
rect 430 10386 99570 10502
rect 9 9494 99600 10386
rect 9 9378 70 9494
rect 430 9378 99570 9494
rect 9 8486 99600 9378
rect 9 8370 70 8486
rect 430 8370 99570 8486
rect 9 7478 99600 8370
rect 9 7362 70 7478
rect 430 7362 99570 7478
rect 9 6806 99600 7362
rect 9 6690 70 6806
rect 430 6690 99570 6806
rect 9 5798 99600 6690
rect 9 5682 70 5798
rect 430 5682 99570 5798
rect 9 4790 99600 5682
rect 9 4674 70 4790
rect 430 4674 99570 4790
rect 9 3782 99600 4674
rect 9 3666 70 3782
rect 430 3666 99570 3782
rect 9 2774 99600 3666
rect 9 2658 70 2774
rect 430 2658 99570 2774
rect 9 1766 99600 2658
rect 9 1650 70 1766
rect 430 1650 99570 1766
rect 9 798 99600 1650
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
<< obsm4 >>
rect 910 32545 2194 55599
rect 2414 32545 9874 55599
rect 10094 32545 17554 55599
rect 17774 32545 17850 55599
<< labels >>
rlabel metal3 s 100 69216 400 69272 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 70224 400 70280 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 34608 400 34664 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 60480 400 60536 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 41328 400 41384 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 35616 400 35672 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 52752 99600 52808 99900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 99600 20160 99900 20216 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 99600 94080 99900 94136 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 67200 99600 67256 99900 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 98112 100 98168 400 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12432 99600 12488 99900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 79632 99600 79688 99900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 70224 100 70280 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 99792 99600 99848 99900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 99600 86352 99900 86408 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 82656 100 82712 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 13440 100 13496 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 83664 400 83720 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 68208 400 68264 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 77952 400 78008 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 62496 400 62552 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 99600 99120 99900 99176 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 65184 100 65240 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 42336 400 42392 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 84672 100 84728 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 10416 400 10472 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 100 89376 400 89432 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 89376 99600 89432 99900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 99600 88368 99900 88424 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 99600 75936 99900 75992 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 99600 98112 99900 98168 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 99600 45024 99900 45080 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 19152 400 19208 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 99600 19152 99900 19208 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 81648 99600 81704 99900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 46032 400 46088 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 51744 400 51800 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 99600 70224 99900 70280 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 99600 64176 99900 64232 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 3696 99600 3752 99900 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 61488 100 61544 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 25872 400 25928 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 91392 100 91448 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 63504 99600 63560 99900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 28560 100 28616 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 9408 100 9464 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 4704 99600 4760 99900 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 35616 99600 35672 99900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 26880 99600 26936 99900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 57456 99600 57512 99900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 85680 100 85736 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 99600 25872 99900 25928 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 97104 99600 97160 99900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 28560 400 28616 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 14112 400 14168 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 100 91392 400 91448 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 83664 100 83720 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 1680 99600 1736 99900 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 99600 50736 99900 50792 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 99600 38304 99900 38360 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 94080 100 94136 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 30576 400 30632 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 87360 99600 87416 99900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 99600 16128 99900 16184 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 81648 400 81704 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 99600 90384 99900 90440 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 55776 99600 55832 99900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 99600 40320 99900 40376 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 74928 400 74984 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 13440 400 13496 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 72912 99600 72968 99900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 78624 400 78680 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 48048 99600 48104 99900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 49728 400 49784 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 99600 97104 99900 97160 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 16128 99600 16184 99900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 30576 99600 30632 99900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 64176 100 64232 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 98112 99600 98168 99900 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 99792 400 99848 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 73920 400 73976 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 40320 100 40376 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 99600 83664 99900 83720 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 11424 100 11480 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 93072 100 93128 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 21840 99600 21896 99900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6720 100 6776 400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 99600 9408 99900 9464 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 66192 400 66248 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 99600 21840 99900 21896 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 37296 400 37352 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 87360 100 87416 400 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 99600 2688 99900 2744 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42336 100 42392 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 33600 100 33656 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 70224 99600 70280 99900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 68208 100 68264 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 99600 35616 99900 35672 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 91392 99600 91448 99900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 35616 100 35672 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 62496 99600 62552 99900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 36288 400 36344 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 66192 100 66248 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 59472 100 59528 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 23856 100 23912 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 4704 400 4760 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 46032 99600 46088 99900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 46032 100 46088 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 42336 99600 42392 99900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 18144 400 18200 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 56784 400 56840 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 72912 100 72968 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 50736 400 50792 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 99600 93072 99900 93128 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 99600 44016 99900 44072 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 30576 100 30632 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 40320 99600 40376 99900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 100 87360 400 87416 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 99600 71904 99900 71960 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 9408 99600 9464 99900 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 99600 15120 99900 15176 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 49728 99600 49784 99900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 15120 400 15176 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 22848 99600 22904 99900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 99600 21168 99900 21224 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 75936 400 75992 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 44016 400 44072 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 99600 74928 99900 74984 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 50736 99600 50792 99900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 21168 99600 21224 99900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 61488 99600 61544 99900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 100 90384 400 90440 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 94080 400 94136 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 99600 24864 99900 24920 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 44016 99600 44072 99900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 7392 400 7448 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 84672 99600 84728 99900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 40320 400 40376 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 67200 400 67256 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 7392 99600 7448 99900 6 la_data_in[34]
port 142 nsew signal input
rlabel metal3 s 100 88368 400 88424 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 71232 100 71288 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal3 s 100 98112 400 98168 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 45024 100 45080 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 54768 99600 54824 99900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 99600 54768 99900 54824 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 34608 100 34664 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 48048 100 48104 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 33600 400 33656 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 94080 99600 94136 99900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 99600 672 99900 728 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 32592 100 32648 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 99600 72912 99900 72968 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 62496 100 62552 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 47040 99600 47096 99900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 38304 99600 38360 99900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 8400 99600 8456 99900 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 39312 99600 39368 99900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 47040 100 47096 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 99600 33600 99900 33656 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 77952 99600 78008 99900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 71232 99600 71288 99900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 26880 400 26936 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 29568 400 29624 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 2688 99600 2744 99900 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 36288 100 36344 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 99600 91392 99900 91448 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 17136 100 17192 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 99600 66192 99900 66248 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 2688 400 2744 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 58464 100 58520 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 25872 99600 25928 99900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 20160 100 20216 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 99600 36288 99900 36344 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1680 400 1736 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 90384 99600 90440 99900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 86352 99600 86408 99900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 99600 53760 99900 53816 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 3696 400 3752 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 71904 400 71960 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 37296 100 37352 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 99600 41328 99900 41384 6 la_data_out[14]
port 184 nsew signal output
rlabel metal3 s 100 85680 400 85736 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 99600 55776 99900 55832 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 49056 99600 49112 99900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 99600 82656 99900 82712 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 52752 100 52808 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 99600 47040 99900 47096 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 99600 14112 99900 14168 6 la_data_out[20]
port 191 nsew signal output
rlabel metal3 s 100 99120 400 99176 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 99600 62496 99900 62552 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 29568 100 29624 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 45024 400 45080 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 53760 100 53816 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 97104 400 97160 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 60480 99600 60536 99900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 99600 79632 99900 79688 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 43008 100 43064 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 22848 400 22904 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 99600 46032 99900 46088 6 la_data_out[30]
port 202 nsew signal output
rlabel metal3 s 99600 4704 99900 4760 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 58464 99600 58520 99900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 99600 18144 99900 18200 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 49056 100 49112 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 53760 99600 53816 99900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 99600 80640 99900 80696 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 99600 39312 99900 39368 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 99600 1680 99900 1736 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 99600 13440 99900 13496 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 16128 400 16184 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 97104 100 97160 400 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 99600 30576 99900 30632 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 99600 84672 99900 84728 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 5712 100 5768 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 41328 100 41384 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 15120 99600 15176 99900 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 14112 99600 14168 99900 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 71232 400 71288 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 22848 100 22904 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 90384 100 90440 400 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 56784 99600 56840 99900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 34608 99600 34664 99900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal3 s 100 96096 400 96152 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 99600 6720 99900 6776 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 95088 400 95144 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 99600 68208 99900 68264 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 37296 99600 37352 99900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 99600 23856 99900 23912 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 75936 99600 75992 99900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 99600 69216 99900 69272 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 38304 400 38360 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 99600 59472 99900 59528 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 80640 99600 80696 99900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 26880 100 26936 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 86352 100 86408 400 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 99600 7392 99900 7448 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 99600 28560 99900 28616 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 96096 99600 96152 99900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 5712 400 5768 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 99600 48048 99900 48104 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 99600 37296 99900 37352 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 99600 71232 99900 71288 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 99600 56784 99900 56840 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 672 99600 728 99900 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 79632 400 79688 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 73920 100 73976 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 88368 100 88424 400 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 14112 100 14168 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 12432 400 12488 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 6720 99600 6776 99900 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 99600 8400 99900 8456 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 19152 99600 19208 99900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 58464 400 58520 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 41328 99600 41384 99900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 73920 99600 73976 99900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 27888 100 27944 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 99600 61488 99900 61544 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 89376 100 89432 400 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 20160 99600 20216 99900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 18144 100 18200 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 61488 400 61544 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 99600 95088 99900 95144 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 99120 99600 99176 99900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 99600 85680 99900 85736 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 43008 99600 43064 99900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 99600 81648 99900 81704 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 50736 100 50792 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 17136 99600 17192 99900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 672 100 728 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 13440 99600 13496 99900 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 51744 100 51800 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 43008 400 43064 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 54768 400 54824 6 la_oenb[3]
port 276 nsew signal input
rlabel metal3 s 99600 12432 99900 12488 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 36288 99600 36344 99900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 63504 400 63560 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 19152 100 19208 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 44016 100 44072 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 82656 99600 82712 99900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 79632 100 79688 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 11424 400 11480 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 72912 400 72968 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 672 400 728 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 100 93072 400 93128 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 76944 100 77000 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 32592 99600 32648 99900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 99120 100 99176 400 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 99600 63504 99900 63560 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 53760 400 53816 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 99600 51744 99900 51800 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 75936 100 75992 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 88368 99600 88424 99900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal3 s 99600 10416 99900 10472 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 59472 99600 59528 99900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 92400 100 92456 400 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 49056 400 49112 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 12432 100 12488 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 99600 50064 99900 50120 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 23856 400 23912 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 99600 65184 99900 65240 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 24864 100 24920 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 95088 100 95144 400 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 28560 99600 28616 99900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 85680 99600 85736 99900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 99600 76944 99900 77000 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 24864 99600 24920 99900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 64176 400 64232 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 99600 17136 99900 17192 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 18144 99600 18200 99900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 99600 34608 99900 34664 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 66192 99600 66248 99900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 45024 99600 45080 99900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 57456 400 57512 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 55776 100 55832 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 9408 400 9464 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 99600 67200 99900 67256 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 63504 100 63560 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 55776 400 55832 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 99600 31584 99900 31640 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 96096 100 96152 400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 93072 99600 93128 99900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 56784 100 56840 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 80640 100 80696 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 99600 22848 99900 22904 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 11424 99600 11480 99900 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 17136 400 17192 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 10416 100 10472 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 33600 99600 33656 99900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 99600 58464 99900 58520 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 99600 96096 99900 96152 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 39312 100 39368 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 99600 42336 99900 42392 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 77952 100 78008 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 76944 99600 77000 99900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 74928 100 74984 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 4704 100 4760 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal3 s 99600 0 99900 56 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 99600 26880 99900 26936 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 31584 99600 31640 99900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 99600 87360 99900 87416 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 76944 400 77000 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal3 s 100 84672 400 84728 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 80640 400 80696 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 3696 100 3752 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 21168 400 21224 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 99600 52752 99900 52808 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 57456 100 57512 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 68208 99600 68264 99900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 92400 99600 92456 99900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 5712 99600 5768 99900 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 15120 100 15176 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 47040 400 47096 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 95088 99600 95144 99900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 59472 400 59528 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 99600 78624 99900 78680 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 99600 32592 99900 32648 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 69216 100 69272 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 83664 99600 83720 99900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 23856 99600 23912 99900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 31584 100 31640 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 99600 60480 99900 60536 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 81648 100 81704 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 99600 29568 99900 29624 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 52752 400 52808 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal3 s 99600 3696 99900 3752 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 16128 100 16184 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 50064 100 50120 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 99600 43008 99900 43064 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 78624 99600 78680 99900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 99600 89376 99900 89432 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal3 s 99600 5712 99900 5768 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 20160 400 20216 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 99600 57456 99900 57512 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1680 100 1736 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 99600 92400 99900 92456 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 74928 99600 74984 99900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal3 s 99600 11424 99900 11480 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 71904 99600 71960 99900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 27888 400 27944 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 31584 400 31640 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 67200 100 67256 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 78624 100 78680 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 48048 400 48104 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal3 s 100 86352 400 86408 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 27888 99600 27944 99900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 32592 400 32648 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 21168 100 21224 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 7392 100 7448 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 51744 99600 51800 99900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 29568 99600 29624 99900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 54768 100 54824 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 69216 99600 69272 99900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 99600 27888 99900 27944 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 65184 400 65240 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 99600 77952 99900 78008 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 21840 100 21896 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 38304 100 38360 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 99600 73920 99900 73976 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 60480 100 60536 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 65184 99600 65240 99900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 64176 99600 64232 99900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal3 s 100 92400 400 92456 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 10416 99600 10472 99900 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 71904 100 71960 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 21840 400 21896 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 82656 400 82712 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 99600 49056 99900 49112 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5897592
string GDS_FILE /home/runner/work/gf180-option23ser/gf180-option23ser/openlane/tiny_user_project/runs/22_12_05_13_56/results/signoff/tiny_user_project.magic.gds
string GDS_START 249392
<< end >>

