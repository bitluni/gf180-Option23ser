module option23serMax (
    input wire [7:0] io_in,
    output reg [7:0] io_out
);
parameter WORD_COUNT = 256;

localparam MSB = WORD_COUNT * 8 - 1;

wire clk = io_in[0];
wire reset = io_in[1];
wire write = io_in[2];
wire din = io_in[3];
wire [3:0] bank = io_in[7:4];

reg [11:0] counter;
reg [MSB: 0] buffer;
reg [8 * 8 * 256 - 1: 0] customChars;

wire writeBuffer = (write && bank == 4'b0000);
wire writeCustom = (write && bank != 4'b0000);
wire shiftBuffer = (counter[2:0] == 3'b111);
wire [10:0] selectedColumn = {buffer[7:0], counter[2:0]};

always@(posedge clk or posedge reset) begin
    if(reset)
        counter <= 3'd0;
    else begin
        if(shiftBuffer && !writeBuffer)
            buffer[MSB:0] <= {buffer[7:0], buffer[MSB:8]};
        if(shiftBuffer && writeBuffer)
            buffer[MSB:0] <= {buffer[7:0], din, buffer[MSB-7:8]};
        if(!shiftBuffer && writeBuffer)
            buffer[MSB:0] <= {din, buffer[MSB:MSB-6], buffer[MSB-8:0]};

        if(write && bank[0])
            customChars[{2'b00,counter}] <= din;
        if(write && bank[1])
            customChars[{2'b01,counter}] <= din;
        if(write && bank[2])
            customChars[{2'b10,counter}] <= din;
        if(write && bank[3])
            customChars[{2'b11,counter}] <= din;
        counter <= counter + 1'd1;
    end
end 

always @ (buffer[7:6] or selectedColumn) begin
if(bank[buffer[7:6]])
    io_out <= customChars[selectedColumn + : 8];
else
    case(selectedColumn)
        11'b00000001000: io_out <= 8'b01111110;
        11'b00000001001: io_out <= 8'b10000001;
        11'b00000001010: io_out <= 8'b10010101;
        11'b00000001011: io_out <= 8'b10110001;
        11'b00000001100: io_out <= 8'b10110001;
        11'b00000001101: io_out <= 8'b10010101;
        11'b00000001110: io_out <= 8'b10000001;
        11'b00000001111: io_out <= 8'b01111110;
        11'b00000010000: io_out <= 8'b01111110;
        11'b00000010001: io_out <= 8'b11111111;
        11'b00000010010: io_out <= 8'b11101011;
        11'b00000010011: io_out <= 8'b11001111;
        11'b00000010100: io_out <= 8'b11001111;
        11'b00000010101: io_out <= 8'b11101011;
        11'b00000010110: io_out <= 8'b11111111;
        11'b00000010111: io_out <= 8'b01111110;
        11'b00000011000: io_out <= 8'b00001110;
        11'b00000011001: io_out <= 8'b00011111;
        11'b00000011010: io_out <= 8'b00111111;
        11'b00000011011: io_out <= 8'b01111110;
        11'b00000011100: io_out <= 8'b00111111;
        11'b00000011101: io_out <= 8'b00011111;
        11'b00000011110: io_out <= 8'b00001110;
        11'b00000100000: io_out <= 8'b00001000;
        11'b00000100001: io_out <= 8'b00011100;
        11'b00000100010: io_out <= 8'b00111110;
        11'b00000100011: io_out <= 8'b01111111;
        11'b00000100100: io_out <= 8'b00111110;
        11'b00000100101: io_out <= 8'b00011100;
        11'b00000100110: io_out <= 8'b00001000;
        11'b00000101000: io_out <= 8'b00111000;
        11'b00000101001: io_out <= 8'b00111010;
        11'b00000101010: io_out <= 8'b10011111;
        11'b00000101011: io_out <= 8'b11111111;
        11'b00000101100: io_out <= 8'b10011111;
        11'b00000101101: io_out <= 8'b00111010;
        11'b00000101110: io_out <= 8'b00111000;
        11'b00000110000: io_out <= 8'b00010000;
        11'b00000110001: io_out <= 8'b00111000;
        11'b00000110010: io_out <= 8'b10111100;
        11'b00000110011: io_out <= 8'b11111111;
        11'b00000110100: io_out <= 8'b10111100;
        11'b00000110101: io_out <= 8'b00111000;
        11'b00000110110: io_out <= 8'b00010000;
        11'b00000111010: io_out <= 8'b00011000;
        11'b00000111011: io_out <= 8'b00111100;
        11'b00000111100: io_out <= 8'b00111100;
        11'b00000111101: io_out <= 8'b00011000;
        11'b00001000000: io_out <= 8'b11111111;
        11'b00001000001: io_out <= 8'b11111111;
        11'b00001000010: io_out <= 8'b11100111;
        11'b00001000011: io_out <= 8'b11000011;
        11'b00001000100: io_out <= 8'b11000011;
        11'b00001000101: io_out <= 8'b11100111;
        11'b00001000110: io_out <= 8'b11111111;
        11'b00001000111: io_out <= 8'b11111111;
        11'b00001001001: io_out <= 8'b00111100;
        11'b00001001010: io_out <= 8'b01100110;
        11'b00001001011: io_out <= 8'b01000010;
        11'b00001001100: io_out <= 8'b01000010;
        11'b00001001101: io_out <= 8'b01100110;
        11'b00001001110: io_out <= 8'b00111100;
        11'b00001010000: io_out <= 8'b11111111;
        11'b00001010001: io_out <= 8'b11000011;
        11'b00001010010: io_out <= 8'b10011001;
        11'b00001010011: io_out <= 8'b10111101;
        11'b00001010100: io_out <= 8'b10111101;
        11'b00001010101: io_out <= 8'b10011001;
        11'b00001010110: io_out <= 8'b11000011;
        11'b00001010111: io_out <= 8'b11111111;
        11'b00001011000: io_out <= 8'b01110000;
        11'b00001011001: io_out <= 8'b10001000;
        11'b00001011010: io_out <= 8'b10001000;
        11'b00001011011: io_out <= 8'b10001000;
        11'b00001011100: io_out <= 8'b10001001;
        11'b00001011101: io_out <= 8'b01111101;
        11'b00001011110: io_out <= 8'b00000011;
        11'b00001011111: io_out <= 8'b00001111;
        11'b00001100001: io_out <= 8'b01001110;
        11'b00001100010: io_out <= 8'b01010001;
        11'b00001100011: io_out <= 8'b11110001;
        11'b00001100100: io_out <= 8'b11110001;
        11'b00001100101: io_out <= 8'b01010001;
        11'b00001100110: io_out <= 8'b01001110;
        11'b00001101000: io_out <= 8'b11000000;
        11'b00001101001: io_out <= 8'b11100000;
        11'b00001101010: io_out <= 8'b01111111;
        11'b00001101011: io_out <= 8'b00000101;
        11'b00001101100: io_out <= 8'b00000101;
        11'b00001101101: io_out <= 8'b00000101;
        11'b00001101110: io_out <= 8'b00000101;
        11'b00001101111: io_out <= 8'b00000111;
        11'b00001110000: io_out <= 8'b11000000;
        11'b00001110001: io_out <= 8'b11100000;
        11'b00001110010: io_out <= 8'b01111111;
        11'b00001110011: io_out <= 8'b00000101;
        11'b00001110100: io_out <= 8'b00000101;
        11'b00001110101: io_out <= 8'b01100101;
        11'b00001110110: io_out <= 8'b01110101;
        11'b00001110111: io_out <= 8'b00111111;
        11'b00001111000: io_out <= 8'b01011010;
        11'b00001111001: io_out <= 8'b01011010;
        11'b00001111010: io_out <= 8'b00111100;
        11'b00001111011: io_out <= 8'b11100111;
        11'b00001111100: io_out <= 8'b11100111;
        11'b00001111101: io_out <= 8'b00111100;
        11'b00001111110: io_out <= 8'b01011010;
        11'b00001111111: io_out <= 8'b01011010;
        11'b00010000000: io_out <= 8'b01111111;
        11'b00010000001: io_out <= 8'b00111110;
        11'b00010000010: io_out <= 8'b00111110;
        11'b00010000011: io_out <= 8'b00011100;
        11'b00010000100: io_out <= 8'b00011100;
        11'b00010000101: io_out <= 8'b00001000;
        11'b00010000110: io_out <= 8'b00001000;
        11'b00010001000: io_out <= 8'b00001000;
        11'b00010001001: io_out <= 8'b00001000;
        11'b00010001010: io_out <= 8'b00011100;
        11'b00010001011: io_out <= 8'b00011100;
        11'b00010001100: io_out <= 8'b00111110;
        11'b00010001101: io_out <= 8'b00111110;
        11'b00010001110: io_out <= 8'b01111111;
        11'b00010010001: io_out <= 8'b00100100;
        11'b00010010010: io_out <= 8'b01100110;
        11'b00010010011: io_out <= 8'b11111111;
        11'b00010010100: io_out <= 8'b11111111;
        11'b00010010101: io_out <= 8'b01100110;
        11'b00010010110: io_out <= 8'b00100100;
        11'b00010011010: io_out <= 8'b01011111;
        11'b00010011101: io_out <= 8'b01011111;
        11'b00010100000: io_out <= 8'b00000110;
        11'b00010100001: io_out <= 8'b00001001;
        11'b00010100010: io_out <= 8'b00001001;
        11'b00010100011: io_out <= 8'b01111111;
        11'b00010100100: io_out <= 8'b00000001;
        11'b00010100101: io_out <= 8'b00000001;
        11'b00010100110: io_out <= 8'b01111111;
        11'b00010100111: io_out <= 8'b00000001;
        11'b00010101000: io_out <= 8'b01000000;
        11'b00010101001: io_out <= 8'b11011010;
        11'b00010101010: io_out <= 8'b10100111;
        11'b00010101011: io_out <= 8'b10100101;
        11'b00010101100: io_out <= 8'b11100101;
        11'b00010101101: io_out <= 8'b01011001;
        11'b00010101110: io_out <= 8'b00000011;
        11'b00010101111: io_out <= 8'b00000010;
        11'b00010110001: io_out <= 8'b01110000;
        11'b00010110010: io_out <= 8'b01110000;
        11'b00010110011: io_out <= 8'b01110000;
        11'b00010110100: io_out <= 8'b01110000;
        11'b00010110101: io_out <= 8'b01110000;
        11'b00010110110: io_out <= 8'b01110000;
        11'b00010111000: io_out <= 8'b10000000;
        11'b00010111001: io_out <= 8'b10010100;
        11'b00010111010: io_out <= 8'b10110110;
        11'b00010111011: io_out <= 8'b11111111;
        11'b00010111100: io_out <= 8'b11111111;
        11'b00010111101: io_out <= 8'b10110110;
        11'b00010111110: io_out <= 8'b10010100;
        11'b00010111111: io_out <= 8'b10000000;
        11'b00011000001: io_out <= 8'b00001100;
        11'b00011000010: io_out <= 8'b00000110;
        11'b00011000011: io_out <= 8'b01111111;
        11'b00011000100: io_out <= 8'b00000110;
        11'b00011000101: io_out <= 8'b00001100;
        11'b00011001001: io_out <= 8'b00011000;
        11'b00011001010: io_out <= 8'b00110000;
        11'b00011001011: io_out <= 8'b01111111;
        11'b00011001100: io_out <= 8'b00110000;
        11'b00011001101: io_out <= 8'b00011000;
        11'b00011010000: io_out <= 8'b00001000;
        11'b00011010001: io_out <= 8'b00001000;
        11'b00011010010: io_out <= 8'b00001000;
        11'b00011010011: io_out <= 8'b00101010;
        11'b00011010100: io_out <= 8'b00111110;
        11'b00011010101: io_out <= 8'b00011100;
        11'b00011010110: io_out <= 8'b00001000;
        11'b00011011000: io_out <= 8'b00001000;
        11'b00011011001: io_out <= 8'b00011100;
        11'b00011011010: io_out <= 8'b00111110;
        11'b00011011011: io_out <= 8'b00101010;
        11'b00011011100: io_out <= 8'b00001000;
        11'b00011011101: io_out <= 8'b00001000;
        11'b00011011110: io_out <= 8'b00001000;
        11'b00011100001: io_out <= 8'b00111100;
        11'b00011100010: io_out <= 8'b00100000;
        11'b00011100011: io_out <= 8'b00100000;
        11'b00011100100: io_out <= 8'b00100000;
        11'b00011100101: io_out <= 8'b00100000;
        11'b00011100110: io_out <= 8'b00100000;
        11'b00011101000: io_out <= 8'b00001000;
        11'b00011101001: io_out <= 8'b00011100;
        11'b00011101010: io_out <= 8'b00111110;
        11'b00011101011: io_out <= 8'b00001000;
        11'b00011101100: io_out <= 8'b00001000;
        11'b00011101101: io_out <= 8'b00111110;
        11'b00011101110: io_out <= 8'b00011100;
        11'b00011101111: io_out <= 8'b00001000;
        11'b00011110000: io_out <= 8'b00110000;
        11'b00011110001: io_out <= 8'b00111000;
        11'b00011110010: io_out <= 8'b00111100;
        11'b00011110011: io_out <= 8'b00111110;
        11'b00011110100: io_out <= 8'b00111100;
        11'b00011110101: io_out <= 8'b00111000;
        11'b00011110110: io_out <= 8'b00110000;
        11'b00011111000: io_out <= 8'b00000110;
        11'b00011111001: io_out <= 8'b00001110;
        11'b00011111010: io_out <= 8'b00011110;
        11'b00011111011: io_out <= 8'b00111110;
        11'b00011111100: io_out <= 8'b00011110;
        11'b00011111101: io_out <= 8'b00001110;
        11'b00011111110: io_out <= 8'b00000110;
        11'b00100001010: io_out <= 8'b00000110;
        11'b00100001011: io_out <= 8'b01011111;
        11'b00100001100: io_out <= 8'b00000110;
        11'b00100010010: io_out <= 8'b00000111;
        11'b00100010101: io_out <= 8'b00000111;
        11'b00100011001: io_out <= 8'b00010100;
        11'b00100011010: io_out <= 8'b01111111;
        11'b00100011011: io_out <= 8'b00010100;
        11'b00100011100: io_out <= 8'b00010100;
        11'b00100011101: io_out <= 8'b01111111;
        11'b00100011110: io_out <= 8'b00010100;
        11'b00100100001: io_out <= 8'b00100100;
        11'b00100100010: io_out <= 8'b00101010;
        11'b00100100011: io_out <= 8'b01101011;
        11'b00100100100: io_out <= 8'b01101011;
        11'b00100100101: io_out <= 8'b00101010;
        11'b00100100110: io_out <= 8'b00010010;
        11'b00100101001: io_out <= 8'b01000110;
        11'b00100101010: io_out <= 8'b00100110;
        11'b00100101011: io_out <= 8'b00010000;
        11'b00100101100: io_out <= 8'b00001000;
        11'b00100101101: io_out <= 8'b01100100;
        11'b00100101110: io_out <= 8'b01100010;
        11'b00100110000: io_out <= 8'b00110000;
        11'b00100110001: io_out <= 8'b01001010;
        11'b00100110010: io_out <= 8'b01000101;
        11'b00100110011: io_out <= 8'b01001101;
        11'b00100110100: io_out <= 8'b00110010;
        11'b00100110101: io_out <= 8'b01001000;
        11'b00100110110: io_out <= 8'b01001000;
        11'b00100111010: io_out <= 8'b00000100;
        11'b00100111011: io_out <= 8'b00000011;
        11'b00101000001: io_out <= 8'b00011100;
        11'b00101000010: io_out <= 8'b00100010;
        11'b00101000011: io_out <= 8'b01000001;
        11'b00101001010: io_out <= 8'b01000001;
        11'b00101001011: io_out <= 8'b00100010;
        11'b00101001100: io_out <= 8'b00011100;
        11'b00101010000: io_out <= 8'b00001000;
        11'b00101010001: io_out <= 8'b00101010;
        11'b00101010010: io_out <= 8'b00011100;
        11'b00101010011: io_out <= 8'b00011100;
        11'b00101010100: io_out <= 8'b00011100;
        11'b00101010101: io_out <= 8'b00101010;
        11'b00101010110: io_out <= 8'b00001000;
        11'b00101011001: io_out <= 8'b00001000;
        11'b00101011010: io_out <= 8'b00001000;
        11'b00101011011: io_out <= 8'b00111110;
        11'b00101011100: io_out <= 8'b00001000;
        11'b00101011101: io_out <= 8'b00001000;
        11'b00101100010: io_out <= 8'b10000000;
        11'b00101100011: io_out <= 8'b01100000;
        11'b00101101001: io_out <= 8'b00001000;
        11'b00101101010: io_out <= 8'b00001000;
        11'b00101101011: io_out <= 8'b00001000;
        11'b00101101100: io_out <= 8'b00001000;
        11'b00101101101: io_out <= 8'b00001000;
        11'b00101101110: io_out <= 8'b00001000;
        11'b00101110011: io_out <= 8'b01100000;
        11'b00101111001: io_out <= 8'b01000000;
        11'b00101111010: io_out <= 8'b00100000;
        11'b00101111011: io_out <= 8'b00010000;
        11'b00101111100: io_out <= 8'b00001000;
        11'b00101111101: io_out <= 8'b00000100;
        11'b00101111110: io_out <= 8'b00000010;
        11'b00110000001: io_out <= 8'b00111110;
        11'b00110000010: io_out <= 8'b01100001;
        11'b00110000011: io_out <= 8'b01010001;
        11'b00110000100: io_out <= 8'b01001001;
        11'b00110000101: io_out <= 8'b01000101;
        11'b00110000110: io_out <= 8'b00111110;
        11'b00110001001: io_out <= 8'b01000100;
        11'b00110001010: io_out <= 8'b01000010;
        11'b00110001011: io_out <= 8'b01111111;
        11'b00110001100: io_out <= 8'b01000000;
        11'b00110001101: io_out <= 8'b01000000;
        11'b00110010001: io_out <= 8'b01100010;
        11'b00110010010: io_out <= 8'b01010001;
        11'b00110010011: io_out <= 8'b01010001;
        11'b00110010100: io_out <= 8'b01001001;
        11'b00110010101: io_out <= 8'b01001001;
        11'b00110010110: io_out <= 8'b01100110;
        11'b00110011001: io_out <= 8'b00100010;
        11'b00110011010: io_out <= 8'b01000001;
        11'b00110011011: io_out <= 8'b01001001;
        11'b00110011100: io_out <= 8'b01001001;
        11'b00110011101: io_out <= 8'b01001001;
        11'b00110011110: io_out <= 8'b00110110;
        11'b00110100000: io_out <= 8'b00010000;
        11'b00110100001: io_out <= 8'b00011000;
        11'b00110100010: io_out <= 8'b00010100;
        11'b00110100011: io_out <= 8'b01010010;
        11'b00110100100: io_out <= 8'b01111111;
        11'b00110100101: io_out <= 8'b01010000;
        11'b00110100110: io_out <= 8'b00010000;
        11'b00110101001: io_out <= 8'b00100111;
        11'b00110101010: io_out <= 8'b01000101;
        11'b00110101011: io_out <= 8'b01000101;
        11'b00110101100: io_out <= 8'b01000101;
        11'b00110101101: io_out <= 8'b01000101;
        11'b00110101110: io_out <= 8'b00111001;
        11'b00110110001: io_out <= 8'b00111100;
        11'b00110110010: io_out <= 8'b01001010;
        11'b00110110011: io_out <= 8'b01001001;
        11'b00110110100: io_out <= 8'b01001001;
        11'b00110110101: io_out <= 8'b01001001;
        11'b00110110110: io_out <= 8'b00110000;
        11'b00110111001: io_out <= 8'b00000011;
        11'b00110111010: io_out <= 8'b00000001;
        11'b00110111011: io_out <= 8'b01110001;
        11'b00110111100: io_out <= 8'b00001001;
        11'b00110111101: io_out <= 8'b00000101;
        11'b00110111110: io_out <= 8'b00000011;
        11'b00111000001: io_out <= 8'b00110110;
        11'b00111000010: io_out <= 8'b01001001;
        11'b00111000011: io_out <= 8'b01001001;
        11'b00111000100: io_out <= 8'b01001001;
        11'b00111000101: io_out <= 8'b01001001;
        11'b00111000110: io_out <= 8'b00110110;
        11'b00111001001: io_out <= 8'b00000110;
        11'b00111001010: io_out <= 8'b01001001;
        11'b00111001011: io_out <= 8'b01001001;
        11'b00111001100: io_out <= 8'b01001001;
        11'b00111001101: io_out <= 8'b00101001;
        11'b00111001110: io_out <= 8'b00011110;
        11'b00111010011: io_out <= 8'b01100110;
        11'b00111011010: io_out <= 8'b10000000;
        11'b00111011011: io_out <= 8'b01100110;
        11'b00111100001: io_out <= 8'b00001000;
        11'b00111100010: io_out <= 8'b00010100;
        11'b00111100011: io_out <= 8'b00100010;
        11'b00111100100: io_out <= 8'b01000001;
        11'b00111101001: io_out <= 8'b00100100;
        11'b00111101010: io_out <= 8'b00100100;
        11'b00111101011: io_out <= 8'b00100100;
        11'b00111101100: io_out <= 8'b00100100;
        11'b00111101101: io_out <= 8'b00100100;
        11'b00111101110: io_out <= 8'b00100100;
        11'b00111110011: io_out <= 8'b01000001;
        11'b00111110100: io_out <= 8'b00100010;
        11'b00111110101: io_out <= 8'b00010100;
        11'b00111110110: io_out <= 8'b00001000;
        11'b00111111001: io_out <= 8'b00000010;
        11'b00111111010: io_out <= 8'b00000001;
        11'b00111111011: io_out <= 8'b00000001;
        11'b00111111100: io_out <= 8'b01010001;
        11'b00111111101: io_out <= 8'b00001001;
        11'b00111111110: io_out <= 8'b00000110;
        11'b01000000001: io_out <= 8'b00111110;
        11'b01000000010: io_out <= 8'b01000001;
        11'b01000000011: io_out <= 8'b01011101;
        11'b01000000100: io_out <= 8'b01010101;
        11'b01000000101: io_out <= 8'b01010101;
        11'b01000000110: io_out <= 8'b00011110;
        11'b01000001001: io_out <= 8'b01111100;
        11'b01000001010: io_out <= 8'b00010010;
        11'b01000001011: io_out <= 8'b00010001;
        11'b01000001100: io_out <= 8'b00010001;
        11'b01000001101: io_out <= 8'b00010010;
        11'b01000001110: io_out <= 8'b01111100;
        11'b01000010001: io_out <= 8'b01000001;
        11'b01000010010: io_out <= 8'b01111111;
        11'b01000010011: io_out <= 8'b01001001;
        11'b01000010100: io_out <= 8'b01001001;
        11'b01000010101: io_out <= 8'b01001001;
        11'b01000010110: io_out <= 8'b00110110;
        11'b01000011001: io_out <= 8'b00011100;
        11'b01000011010: io_out <= 8'b00100010;
        11'b01000011011: io_out <= 8'b01000001;
        11'b01000011100: io_out <= 8'b01000001;
        11'b01000011101: io_out <= 8'b01000001;
        11'b01000011110: io_out <= 8'b00100010;
        11'b01000100001: io_out <= 8'b01000001;
        11'b01000100010: io_out <= 8'b01111111;
        11'b01000100011: io_out <= 8'b01000001;
        11'b01000100100: io_out <= 8'b01000001;
        11'b01000100101: io_out <= 8'b00100010;
        11'b01000100110: io_out <= 8'b00011100;
        11'b01000101001: io_out <= 8'b01000001;
        11'b01000101010: io_out <= 8'b01111111;
        11'b01000101011: io_out <= 8'b01001001;
        11'b01000101100: io_out <= 8'b01011101;
        11'b01000101101: io_out <= 8'b01000001;
        11'b01000101110: io_out <= 8'b01100011;
        11'b01000110001: io_out <= 8'b01000001;
        11'b01000110010: io_out <= 8'b01111111;
        11'b01000110011: io_out <= 8'b01001001;
        11'b01000110100: io_out <= 8'b00011101;
        11'b01000110101: io_out <= 8'b00000001;
        11'b01000110110: io_out <= 8'b00000011;
        11'b01000111001: io_out <= 8'b00011100;
        11'b01000111010: io_out <= 8'b00100010;
        11'b01000111011: io_out <= 8'b01000001;
        11'b01000111100: io_out <= 8'b01010001;
        11'b01000111101: io_out <= 8'b01010001;
        11'b01000111110: io_out <= 8'b01110010;
        11'b01001000001: io_out <= 8'b01111111;
        11'b01001000010: io_out <= 8'b00001000;
        11'b01001000011: io_out <= 8'b00001000;
        11'b01001000100: io_out <= 8'b00001000;
        11'b01001000101: io_out <= 8'b00001000;
        11'b01001000110: io_out <= 8'b01111111;
        11'b01001001010: io_out <= 8'b01000001;
        11'b01001001011: io_out <= 8'b01111111;
        11'b01001001100: io_out <= 8'b01000001;
        11'b01001010001: io_out <= 8'b00110000;
        11'b01001010010: io_out <= 8'b01000000;
        11'b01001010011: io_out <= 8'b01000000;
        11'b01001010100: io_out <= 8'b01000001;
        11'b01001010101: io_out <= 8'b00111111;
        11'b01001010110: io_out <= 8'b00000001;
        11'b01001011001: io_out <= 8'b01000001;
        11'b01001011010: io_out <= 8'b01111111;
        11'b01001011011: io_out <= 8'b00001000;
        11'b01001011100: io_out <= 8'b00010100;
        11'b01001011101: io_out <= 8'b00100010;
        11'b01001011110: io_out <= 8'b01000001;
        11'b01001011111: io_out <= 8'b01000000;
        11'b01001100001: io_out <= 8'b01000001;
        11'b01001100010: io_out <= 8'b01111111;
        11'b01001100011: io_out <= 8'b01000001;
        11'b01001100100: io_out <= 8'b01000000;
        11'b01001100101: io_out <= 8'b01000000;
        11'b01001100110: io_out <= 8'b01100000;
        11'b01001101001: io_out <= 8'b01111111;
        11'b01001101010: io_out <= 8'b00000001;
        11'b01001101011: io_out <= 8'b00000010;
        11'b01001101100: io_out <= 8'b00000100;
        11'b01001101101: io_out <= 8'b00000010;
        11'b01001101110: io_out <= 8'b00000001;
        11'b01001101111: io_out <= 8'b01111111;
        11'b01001110001: io_out <= 8'b01111111;
        11'b01001110010: io_out <= 8'b00000001;
        11'b01001110011: io_out <= 8'b00000010;
        11'b01001110100: io_out <= 8'b00000100;
        11'b01001110101: io_out <= 8'b00001000;
        11'b01001110110: io_out <= 8'b01111111;
        11'b01001111001: io_out <= 8'b00011100;
        11'b01001111010: io_out <= 8'b00100010;
        11'b01001111011: io_out <= 8'b01000001;
        11'b01001111100: io_out <= 8'b01000001;
        11'b01001111101: io_out <= 8'b00100010;
        11'b01001111110: io_out <= 8'b00011100;
        11'b01010000001: io_out <= 8'b01000001;
        11'b01010000010: io_out <= 8'b01111111;
        11'b01010000011: io_out <= 8'b01001001;
        11'b01010000100: io_out <= 8'b00001001;
        11'b01010000101: io_out <= 8'b00001001;
        11'b01010000110: io_out <= 8'b00000110;
        11'b01010001001: io_out <= 8'b00011110;
        11'b01010001010: io_out <= 8'b00100001;
        11'b01010001011: io_out <= 8'b00100001;
        11'b01010001100: io_out <= 8'b00110001;
        11'b01010001101: io_out <= 8'b00100001;
        11'b01010001110: io_out <= 8'b01011110;
        11'b01010001111: io_out <= 8'b01000000;
        11'b01010010001: io_out <= 8'b01000001;
        11'b01010010010: io_out <= 8'b01111111;
        11'b01010010011: io_out <= 8'b01001001;
        11'b01010010100: io_out <= 8'b00011001;
        11'b01010010101: io_out <= 8'b00101001;
        11'b01010010110: io_out <= 8'b01000110;
        11'b01010011001: io_out <= 8'b00100110;
        11'b01010011010: io_out <= 8'b01001001;
        11'b01010011011: io_out <= 8'b01001001;
        11'b01010011100: io_out <= 8'b01001001;
        11'b01010011101: io_out <= 8'b01001001;
        11'b01010011110: io_out <= 8'b00110010;
        11'b01010100001: io_out <= 8'b00000011;
        11'b01010100010: io_out <= 8'b00000001;
        11'b01010100011: io_out <= 8'b01000001;
        11'b01010100100: io_out <= 8'b01111111;
        11'b01010100101: io_out <= 8'b01000001;
        11'b01010100110: io_out <= 8'b00000001;
        11'b01010100111: io_out <= 8'b00000011;
        11'b01010101001: io_out <= 8'b00111111;
        11'b01010101010: io_out <= 8'b01000000;
        11'b01010101011: io_out <= 8'b01000000;
        11'b01010101100: io_out <= 8'b01000000;
        11'b01010101101: io_out <= 8'b01000000;
        11'b01010101110: io_out <= 8'b00111111;
        11'b01010110001: io_out <= 8'b00001111;
        11'b01010110010: io_out <= 8'b00010000;
        11'b01010110011: io_out <= 8'b00100000;
        11'b01010110100: io_out <= 8'b01000000;
        11'b01010110101: io_out <= 8'b00100000;
        11'b01010110110: io_out <= 8'b00010000;
        11'b01010110111: io_out <= 8'b00001111;
        11'b01010111001: io_out <= 8'b00111111;
        11'b01010111010: io_out <= 8'b01000000;
        11'b01010111011: io_out <= 8'b01000000;
        11'b01010111100: io_out <= 8'b00111000;
        11'b01010111101: io_out <= 8'b01000000;
        11'b01010111110: io_out <= 8'b01000000;
        11'b01010111111: io_out <= 8'b00111111;
        11'b01011000001: io_out <= 8'b01000001;
        11'b01011000010: io_out <= 8'b00100010;
        11'b01011000011: io_out <= 8'b00010100;
        11'b01011000100: io_out <= 8'b00001000;
        11'b01011000101: io_out <= 8'b00010100;
        11'b01011000110: io_out <= 8'b00100010;
        11'b01011000111: io_out <= 8'b01000001;
        11'b01011001001: io_out <= 8'b00000001;
        11'b01011001010: io_out <= 8'b00000010;
        11'b01011001011: io_out <= 8'b01000100;
        11'b01011001100: io_out <= 8'b01111000;
        11'b01011001101: io_out <= 8'b01000100;
        11'b01011001110: io_out <= 8'b00000010;
        11'b01011001111: io_out <= 8'b00000001;
        11'b01011010001: io_out <= 8'b01000011;
        11'b01011010010: io_out <= 8'b01100001;
        11'b01011010011: io_out <= 8'b01010001;
        11'b01011010100: io_out <= 8'b01001001;
        11'b01011010101: io_out <= 8'b01000101;
        11'b01011010110: io_out <= 8'b01000011;
        11'b01011010111: io_out <= 8'b01100001;
        11'b01011011001: io_out <= 8'b01111111;
        11'b01011011010: io_out <= 8'b01000001;
        11'b01011011011: io_out <= 8'b01000001;
        11'b01011011100: io_out <= 8'b01000001;
        11'b01011100000: io_out <= 8'b00000001;
        11'b01011100001: io_out <= 8'b00000010;
        11'b01011100010: io_out <= 8'b00000100;
        11'b01011100011: io_out <= 8'b00001000;
        11'b01011100100: io_out <= 8'b00010000;
        11'b01011100101: io_out <= 8'b00100000;
        11'b01011100110: io_out <= 8'b01000000;
        11'b01011101001: io_out <= 8'b01000001;
        11'b01011101010: io_out <= 8'b01000001;
        11'b01011101011: io_out <= 8'b01000001;
        11'b01011101100: io_out <= 8'b01111111;
        11'b01011110000: io_out <= 8'b00001000;
        11'b01011110001: io_out <= 8'b00000100;
        11'b01011110010: io_out <= 8'b00000010;
        11'b01011110011: io_out <= 8'b00000001;
        11'b01011110100: io_out <= 8'b00000010;
        11'b01011110101: io_out <= 8'b00000100;
        11'b01011110110: io_out <= 8'b00001000;
        11'b01011111000: io_out <= 8'b10000000;
        11'b01011111001: io_out <= 8'b10000000;
        11'b01011111010: io_out <= 8'b10000000;
        11'b01011111011: io_out <= 8'b10000000;
        11'b01011111100: io_out <= 8'b10000000;
        11'b01011111101: io_out <= 8'b10000000;
        11'b01011111110: io_out <= 8'b10000000;
        11'b01011111111: io_out <= 8'b10000000;
        11'b01100000011: io_out <= 8'b00000011;
        11'b01100000100: io_out <= 8'b00000100;
        11'b01100001001: io_out <= 8'b00100000;
        11'b01100001010: io_out <= 8'b01010100;
        11'b01100001011: io_out <= 8'b01010100;
        11'b01100001100: io_out <= 8'b01010100;
        11'b01100001101: io_out <= 8'b01010100;
        11'b01100001110: io_out <= 8'b01111000;
        11'b01100001111: io_out <= 8'b01000000;
        11'b01100010001: io_out <= 8'b00000001;
        11'b01100010010: io_out <= 8'b01111111;
        11'b01100010011: io_out <= 8'b00110000;
        11'b01100010100: io_out <= 8'b01001000;
        11'b01100010101: io_out <= 8'b01001000;
        11'b01100010110: io_out <= 8'b01001000;
        11'b01100010111: io_out <= 8'b00110000;
        11'b01100011001: io_out <= 8'b00111000;
        11'b01100011010: io_out <= 8'b01000100;
        11'b01100011011: io_out <= 8'b01000100;
        11'b01100011100: io_out <= 8'b01000100;
        11'b01100011101: io_out <= 8'b01000100;
        11'b01100011110: io_out <= 8'b00101000;
        11'b01100100001: io_out <= 8'b00110000;
        11'b01100100010: io_out <= 8'b01001000;
        11'b01100100011: io_out <= 8'b01001000;
        11'b01100100100: io_out <= 8'b01001000;
        11'b01100100101: io_out <= 8'b00110001;
        11'b01100100110: io_out <= 8'b01111111;
        11'b01100100111: io_out <= 8'b01000000;
        11'b01100101001: io_out <= 8'b00111000;
        11'b01100101010: io_out <= 8'b01010100;
        11'b01100101011: io_out <= 8'b01010100;
        11'b01100101100: io_out <= 8'b01010100;
        11'b01100101101: io_out <= 8'b01010100;
        11'b01100101110: io_out <= 8'b00011000;
        11'b01100110010: io_out <= 8'b01001000;
        11'b01100110011: io_out <= 8'b01111110;
        11'b01100110100: io_out <= 8'b01001001;
        11'b01100110101: io_out <= 8'b00000001;
        11'b01100110110: io_out <= 8'b00000010;
        11'b01100111001: io_out <= 8'b10011000;
        11'b01100111010: io_out <= 8'b10100100;
        11'b01100111011: io_out <= 8'b10100100;
        11'b01100111100: io_out <= 8'b10100100;
        11'b01100111101: io_out <= 8'b10100100;
        11'b01100111110: io_out <= 8'b01111000;
        11'b01100111111: io_out <= 8'b00000100;
        11'b01101000001: io_out <= 8'b01000001;
        11'b01101000010: io_out <= 8'b01111111;
        11'b01101000011: io_out <= 8'b00001000;
        11'b01101000100: io_out <= 8'b00000100;
        11'b01101000101: io_out <= 8'b00000100;
        11'b01101000110: io_out <= 8'b01111000;
        11'b01101001010: io_out <= 8'b01000100;
        11'b01101001011: io_out <= 8'b01111101;
        11'b01101001100: io_out <= 8'b01000000;
        11'b01101010001: io_out <= 8'b01100000;
        11'b01101010010: io_out <= 8'b10000000;
        11'b01101010011: io_out <= 8'b10000000;
        11'b01101010100: io_out <= 8'b10000000;
        11'b01101010101: io_out <= 8'b10000100;
        11'b01101010110: io_out <= 8'b01111101;
        11'b01101011001: io_out <= 8'b00000001;
        11'b01101011010: io_out <= 8'b01111111;
        11'b01101011011: io_out <= 8'b00010000;
        11'b01101011100: io_out <= 8'b00101000;
        11'b01101011101: io_out <= 8'b01000100;
        11'b01101011110: io_out <= 8'b01000000;
        11'b01101100010: io_out <= 8'b01000001;
        11'b01101100011: io_out <= 8'b01111111;
        11'b01101100100: io_out <= 8'b01000000;
        11'b01101101001: io_out <= 8'b01111100;
        11'b01101101010: io_out <= 8'b00000100;
        11'b01101101011: io_out <= 8'b00000100;
        11'b01101101100: io_out <= 8'b01111000;
        11'b01101101101: io_out <= 8'b00000100;
        11'b01101101110: io_out <= 8'b00000100;
        11'b01101101111: io_out <= 8'b01111000;
        11'b01101110001: io_out <= 8'b01111100;
        11'b01101110010: io_out <= 8'b00001000;
        11'b01101110011: io_out <= 8'b00000100;
        11'b01101110100: io_out <= 8'b00000100;
        11'b01101110101: io_out <= 8'b00000100;
        11'b01101110110: io_out <= 8'b01111000;
        11'b01101111001: io_out <= 8'b00111000;
        11'b01101111010: io_out <= 8'b01000100;
        11'b01101111011: io_out <= 8'b01000100;
        11'b01101111100: io_out <= 8'b01000100;
        11'b01101111101: io_out <= 8'b01000100;
        11'b01101111110: io_out <= 8'b00111000;
        11'b01110000001: io_out <= 8'b10000100;
        11'b01110000010: io_out <= 8'b11111100;
        11'b01110000011: io_out <= 8'b10011000;
        11'b01110000100: io_out <= 8'b00100100;
        11'b01110000101: io_out <= 8'b00100100;
        11'b01110000110: io_out <= 8'b00011000;
        11'b01110001001: io_out <= 8'b00011000;
        11'b01110001010: io_out <= 8'b00100100;
        11'b01110001011: io_out <= 8'b00100100;
        11'b01110001100: io_out <= 8'b10011000;
        11'b01110001101: io_out <= 8'b11111100;
        11'b01110001110: io_out <= 8'b10000100;
        11'b01110010001: io_out <= 8'b01000100;
        11'b01110010010: io_out <= 8'b01111100;
        11'b01110010011: io_out <= 8'b01001000;
        11'b01110010100: io_out <= 8'b00000100;
        11'b01110010101: io_out <= 8'b00000100;
        11'b01110010110: io_out <= 8'b00011000;
        11'b01110011001: io_out <= 8'b01001000;
        11'b01110011010: io_out <= 8'b01010100;
        11'b01110011011: io_out <= 8'b01010100;
        11'b01110011100: io_out <= 8'b01010100;
        11'b01110011101: io_out <= 8'b01010100;
        11'b01110011110: io_out <= 8'b00100100;
        11'b01110100001: io_out <= 8'b00000100;
        11'b01110100010: io_out <= 8'b00000100;
        11'b01110100011: io_out <= 8'b00111111;
        11'b01110100100: io_out <= 8'b01000100;
        11'b01110100101: io_out <= 8'b01000100;
        11'b01110100110: io_out <= 8'b00100000;
        11'b01110101001: io_out <= 8'b00111100;
        11'b01110101010: io_out <= 8'b01000000;
        11'b01110101011: io_out <= 8'b01000000;
        11'b01110101100: io_out <= 8'b01000000;
        11'b01110101101: io_out <= 8'b00100000;
        11'b01110101110: io_out <= 8'b01111100;
        11'b01110110001: io_out <= 8'b00001100;
        11'b01110110010: io_out <= 8'b00010000;
        11'b01110110011: io_out <= 8'b00100000;
        11'b01110110100: io_out <= 8'b01000000;
        11'b01110110101: io_out <= 8'b00100000;
        11'b01110110110: io_out <= 8'b00010000;
        11'b01110110111: io_out <= 8'b00001100;
        11'b01110111001: io_out <= 8'b00111100;
        11'b01110111010: io_out <= 8'b01000000;
        11'b01110111011: io_out <= 8'b01000000;
        11'b01110111100: io_out <= 8'b00111000;
        11'b01110111101: io_out <= 8'b01000000;
        11'b01110111110: io_out <= 8'b01000000;
        11'b01110111111: io_out <= 8'b00111100;
        11'b01111000001: io_out <= 8'b01000100;
        11'b01111000010: io_out <= 8'b00101000;
        11'b01111000011: io_out <= 8'b00010000;
        11'b01111000100: io_out <= 8'b00101000;
        11'b01111000101: io_out <= 8'b01000100;
        11'b01111001001: io_out <= 8'b10011100;
        11'b01111001010: io_out <= 8'b10100000;
        11'b01111001011: io_out <= 8'b10100000;
        11'b01111001100: io_out <= 8'b10100000;
        11'b01111001101: io_out <= 8'b10100000;
        11'b01111001110: io_out <= 8'b01111100;
        11'b01111010001: io_out <= 8'b01000100;
        11'b01111010010: io_out <= 8'b01100100;
        11'b01111010011: io_out <= 8'b01010100;
        11'b01111010100: io_out <= 8'b01001100;
        11'b01111010101: io_out <= 8'b01000100;
        11'b01111011001: io_out <= 8'b00001000;
        11'b01111011010: io_out <= 8'b00001000;
        11'b01111011011: io_out <= 8'b00110110;
        11'b01111011100: io_out <= 8'b01000001;
        11'b01111011101: io_out <= 8'b01000001;
        11'b01111100011: io_out <= 8'b01110111;
        11'b01111101010: io_out <= 8'b01000001;
        11'b01111101011: io_out <= 8'b01000001;
        11'b01111101100: io_out <= 8'b00110110;
        11'b01111101101: io_out <= 8'b00001000;
        11'b01111101110: io_out <= 8'b00001000;
        11'b01111110001: io_out <= 8'b00000010;
        11'b01111110010: io_out <= 8'b00000001;
        11'b01111110011: io_out <= 8'b00000001;
        11'b01111110100: io_out <= 8'b00000010;
        11'b01111110101: io_out <= 8'b00000010;
        11'b01111110110: io_out <= 8'b00000001;
        11'b01111111001: io_out <= 8'b01110000;
        11'b01111111010: io_out <= 8'b01001000;
        11'b01111111011: io_out <= 8'b01000100;
        11'b01111111100: io_out <= 8'b01000010;
        11'b01111111101: io_out <= 8'b01000100;
        11'b01111111110: io_out <= 8'b01001000;
        11'b01111111111: io_out <= 8'b01110000;
        11'b10000000001: io_out <= 8'b00001110;
        11'b10000000010: io_out <= 8'b10010001;
        11'b10000000011: io_out <= 8'b10010001;
        11'b10000000100: io_out <= 8'b10110001;
        11'b10000000101: io_out <= 8'b10110001;
        11'b10000000110: io_out <= 8'b01001010;
        11'b10000001001: io_out <= 8'b00111010;
        11'b10000001010: io_out <= 8'b01000000;
        11'b10000001011: io_out <= 8'b01000000;
        11'b10000001100: io_out <= 8'b01000000;
        11'b10000001101: io_out <= 8'b01111010;
        11'b10000001110: io_out <= 8'b01000000;
        11'b10000010001: io_out <= 8'b00111000;
        11'b10000010010: io_out <= 8'b01010100;
        11'b10000010011: io_out <= 8'b01010100;
        11'b10000010100: io_out <= 8'b01010101;
        11'b10000010101: io_out <= 8'b01010101;
        11'b10000010110: io_out <= 8'b00011000;
        11'b10000011001: io_out <= 8'b00100010;
        11'b10000011010: io_out <= 8'b01010101;
        11'b10000011011: io_out <= 8'b01010101;
        11'b10000011100: io_out <= 8'b01010101;
        11'b10000011101: io_out <= 8'b01111001;
        11'b10000011110: io_out <= 8'b01000010;
        11'b10000100001: io_out <= 8'b00100001;
        11'b10000100010: io_out <= 8'b01010100;
        11'b10000100011: io_out <= 8'b01010100;
        11'b10000100100: io_out <= 8'b01010100;
        11'b10000100101: io_out <= 8'b01111000;
        11'b10000100110: io_out <= 8'b01000001;
        11'b10000101001: io_out <= 8'b00100000;
        11'b10000101010: io_out <= 8'b01010101;
        11'b10000101011: io_out <= 8'b01010101;
        11'b10000101100: io_out <= 8'b01010100;
        11'b10000101101: io_out <= 8'b01111000;
        11'b10000101110: io_out <= 8'b01000000;
        11'b10000110001: io_out <= 8'b00100000;
        11'b10000110010: io_out <= 8'b01010100;
        11'b10000110011: io_out <= 8'b01010101;
        11'b10000110100: io_out <= 8'b01010100;
        11'b10000110101: io_out <= 8'b01111000;
        11'b10000110110: io_out <= 8'b01000000;
        11'b10000111001: io_out <= 8'b00011000;
        11'b10000111010: io_out <= 8'b00100100;
        11'b10000111011: io_out <= 8'b10100100;
        11'b10000111100: io_out <= 8'b10100100;
        11'b10000111101: io_out <= 8'b11100100;
        11'b10000111110: io_out <= 8'b01000000;
        11'b10001000001: io_out <= 8'b00111010;
        11'b10001000010: io_out <= 8'b01010101;
        11'b10001000011: io_out <= 8'b01010101;
        11'b10001000100: io_out <= 8'b01010101;
        11'b10001000101: io_out <= 8'b01010101;
        11'b10001000110: io_out <= 8'b00011010;
        11'b10001001001: io_out <= 8'b00111001;
        11'b10001001010: io_out <= 8'b01010100;
        11'b10001001011: io_out <= 8'b01010100;
        11'b10001001100: io_out <= 8'b01010100;
        11'b10001001101: io_out <= 8'b01010100;
        11'b10001001110: io_out <= 8'b00011001;
        11'b10001010001: io_out <= 8'b00111000;
        11'b10001010010: io_out <= 8'b01010101;
        11'b10001010011: io_out <= 8'b01010101;
        11'b10001010100: io_out <= 8'b01010100;
        11'b10001010101: io_out <= 8'b01010100;
        11'b10001010110: io_out <= 8'b00011000;
        11'b10001011010: io_out <= 8'b00000001;
        11'b10001011011: io_out <= 8'b01000100;
        11'b10001011100: io_out <= 8'b01111100;
        11'b10001011101: io_out <= 8'b01000001;
        11'b10001100000: io_out <= 8'b00000010;
        11'b10001100001: io_out <= 8'b00000001;
        11'b10001100010: io_out <= 8'b01000101;
        11'b10001100011: io_out <= 8'b01111101;
        11'b10001100100: io_out <= 8'b01000001;
        11'b10001100101: io_out <= 8'b00000001;
        11'b10001100110: io_out <= 8'b00000010;
        11'b10001101010: io_out <= 8'b00000001;
        11'b10001101011: io_out <= 8'b01000101;
        11'b10001101100: io_out <= 8'b01111100;
        11'b10001101101: io_out <= 8'b01000000;
        11'b10001110001: io_out <= 8'b01111001;
        11'b10001110010: io_out <= 8'b00010100;
        11'b10001110011: io_out <= 8'b00010010;
        11'b10001110100: io_out <= 8'b00010010;
        11'b10001110101: io_out <= 8'b00010100;
        11'b10001110110: io_out <= 8'b01111001;
        11'b10001111001: io_out <= 8'b01110000;
        11'b10001111010: io_out <= 8'b00101000;
        11'b10001111011: io_out <= 8'b00101011;
        11'b10001111100: io_out <= 8'b00101011;
        11'b10001111101: io_out <= 8'b00101000;
        11'b10001111110: io_out <= 8'b01110000;
        11'b10010000001: io_out <= 8'b01000100;
        11'b10010000010: io_out <= 8'b01111100;
        11'b10010000011: io_out <= 8'b01010100;
        11'b10010000100: io_out <= 8'b01010101;
        11'b10010000101: io_out <= 8'b01000101;
        11'b10010001001: io_out <= 8'b00100000;
        11'b10010001010: io_out <= 8'b01010100;
        11'b10010001011: io_out <= 8'b01010100;
        11'b10010001100: io_out <= 8'b01011000;
        11'b10010001101: io_out <= 8'b00111000;
        11'b10010001110: io_out <= 8'b01010100;
        11'b10010001111: io_out <= 8'b01010100;
        11'b10010010001: io_out <= 8'b01111100;
        11'b10010010010: io_out <= 8'b00001010;
        11'b10010010011: io_out <= 8'b00001001;
        11'b10010010100: io_out <= 8'b00001001;
        11'b10010010101: io_out <= 8'b01111111;
        11'b10010010110: io_out <= 8'b01001001;
        11'b10010010111: io_out <= 8'b01001001;
        11'b10010011001: io_out <= 8'b00110000;
        11'b10010011010: io_out <= 8'b01001010;
        11'b10010011011: io_out <= 8'b01001001;
        11'b10010011100: io_out <= 8'b01001001;
        11'b10010011101: io_out <= 8'b01001010;
        11'b10010011110: io_out <= 8'b00110000;
        11'b10010100001: io_out <= 8'b00110010;
        11'b10010100010: io_out <= 8'b01001000;
        11'b10010100011: io_out <= 8'b01001000;
        11'b10010100100: io_out <= 8'b01001000;
        11'b10010100101: io_out <= 8'b01001000;
        11'b10010100110: io_out <= 8'b00110010;
        11'b10010101001: io_out <= 8'b00110000;
        11'b10010101010: io_out <= 8'b01001001;
        11'b10010101011: io_out <= 8'b01001010;
        11'b10010101100: io_out <= 8'b01001000;
        11'b10010101101: io_out <= 8'b01001000;
        11'b10010101110: io_out <= 8'b00110000;
        11'b10010110001: io_out <= 8'b00111000;
        11'b10010110010: io_out <= 8'b01000010;
        11'b10010110011: io_out <= 8'b01000001;
        11'b10010110100: io_out <= 8'b01000001;
        11'b10010110101: io_out <= 8'b01000010;
        11'b10010110110: io_out <= 8'b00111000;
        11'b10010111001: io_out <= 8'b00111000;
        11'b10010111010: io_out <= 8'b01000001;
        11'b10010111011: io_out <= 8'b01000010;
        11'b10010111100: io_out <= 8'b01000000;
        11'b10010111101: io_out <= 8'b01000000;
        11'b10010111110: io_out <= 8'b00111000;
        11'b10011000001: io_out <= 8'b00011010;
        11'b10011000010: io_out <= 8'b10100000;
        11'b10011000011: io_out <= 8'b10100000;
        11'b10011000100: io_out <= 8'b10100000;
        11'b10011000101: io_out <= 8'b10100000;
        11'b10011000110: io_out <= 8'b01111010;
        11'b10011001001: io_out <= 8'b00011001;
        11'b10011001010: io_out <= 8'b00100100;
        11'b10011001011: io_out <= 8'b01000010;
        11'b10011001100: io_out <= 8'b01000010;
        11'b10011001101: io_out <= 8'b00100100;
        11'b10011001110: io_out <= 8'b00011001;
        11'b10011010001: io_out <= 8'b00111101;
        11'b10011010010: io_out <= 8'b01000000;
        11'b10011010011: io_out <= 8'b01000000;
        11'b10011010100: io_out <= 8'b01000000;
        11'b10011010101: io_out <= 8'b01000000;
        11'b10011010110: io_out <= 8'b00111101;
        11'b10011011001: io_out <= 8'b00011000;
        11'b10011011010: io_out <= 8'b00100100;
        11'b10011011011: io_out <= 8'b00100100;
        11'b10011011100: io_out <= 8'b11100111;
        11'b10011011101: io_out <= 8'b00100100;
        11'b10011011110: io_out <= 8'b00100100;
        11'b10011100001: io_out <= 8'b01101000;
        11'b10011100010: io_out <= 8'b01011110;
        11'b10011100011: io_out <= 8'b01001001;
        11'b10011100100: io_out <= 8'b01000001;
        11'b10011100101: io_out <= 8'b01000010;
        11'b10011100110: io_out <= 8'b00100000;
        11'b10011101001: io_out <= 8'b00010101;
        11'b10011101010: io_out <= 8'b00010110;
        11'b10011101011: io_out <= 8'b01111100;
        11'b10011101100: io_out <= 8'b00010110;
        11'b10011101101: io_out <= 8'b00010101;
        11'b10011110000: io_out <= 8'b10000001;
        11'b10011110001: io_out <= 8'b11111111;
        11'b10011110010: io_out <= 8'b10000101;
        11'b10011110011: io_out <= 8'b00000101;
        11'b10011110100: io_out <= 8'b00010111;
        11'b10011110101: io_out <= 8'b11111010;
        11'b10011110110: io_out <= 8'b10010000;
        11'b10011110111: io_out <= 8'b01010000;
        11'b10011111000: io_out <= 8'b01000000;
        11'b10011111001: io_out <= 8'b10001000;
        11'b10011111010: io_out <= 8'b10001000;
        11'b10011111011: io_out <= 8'b01111111;
        11'b10011111100: io_out <= 8'b00001001;
        11'b10011111101: io_out <= 8'b00001001;
        11'b10011111110: io_out <= 8'b00000010;
        11'b10100000001: io_out <= 8'b00100000;
        11'b10100000010: io_out <= 8'b01010100;
        11'b10100000011: io_out <= 8'b01010100;
        11'b10100000100: io_out <= 8'b01010101;
        11'b10100000101: io_out <= 8'b01111001;
        11'b10100000110: io_out <= 8'b01000000;
        11'b10100001011: io_out <= 8'b01000100;
        11'b10100001100: io_out <= 8'b01111101;
        11'b10100001101: io_out <= 8'b01000001;
        11'b10100010001: io_out <= 8'b00110000;
        11'b10100010010: io_out <= 8'b01001000;
        11'b10100010011: io_out <= 8'b01001000;
        11'b10100010100: io_out <= 8'b01001010;
        11'b10100010101: io_out <= 8'b01001001;
        11'b10100010110: io_out <= 8'b00110000;
        11'b10100011001: io_out <= 8'b00111000;
        11'b10100011010: io_out <= 8'b01000000;
        11'b10100011011: io_out <= 8'b01000000;
        11'b10100011100: io_out <= 8'b01000100;
        11'b10100011101: io_out <= 8'b01000010;
        11'b10100011110: io_out <= 8'b00111000;
        11'b10100100001: io_out <= 8'b01111010;
        11'b10100100010: io_out <= 8'b00001001;
        11'b10100100011: io_out <= 8'b00001001;
        11'b10100100100: io_out <= 8'b00001010;
        11'b10100100101: io_out <= 8'b00001010;
        11'b10100100110: io_out <= 8'b01110001;
        11'b10100101001: io_out <= 8'b01111010;
        11'b10100101010: io_out <= 8'b00001001;
        11'b10100101011: io_out <= 8'b00010001;
        11'b10100101100: io_out <= 8'b00100010;
        11'b10100101101: io_out <= 8'b01000011;
        11'b10100101110: io_out <= 8'b01111000;
        11'b10100110001: io_out <= 8'b00100110;
        11'b10100110010: io_out <= 8'b00101001;
        11'b10100110011: io_out <= 8'b00101001;
        11'b10100110100: io_out <= 8'b00101001;
        11'b10100110101: io_out <= 8'b00101111;
        11'b10100110110: io_out <= 8'b00101000;
        11'b10100111001: io_out <= 8'b00100110;
        11'b10100111010: io_out <= 8'b00101001;
        11'b10100111011: io_out <= 8'b00101001;
        11'b10100111100: io_out <= 8'b00101001;
        11'b10100111101: io_out <= 8'b00100110;
        11'b10101000001: io_out <= 8'b00110000;
        11'b10101000010: io_out <= 8'b01001000;
        11'b10101000011: io_out <= 8'b01000101;
        11'b10101000100: io_out <= 8'b01000000;
        11'b10101000101: io_out <= 8'b01000000;
        11'b10101000110: io_out <= 8'b00100000;
        11'b10101001001: io_out <= 8'b00111000;
        11'b10101001010: io_out <= 8'b00001000;
        11'b10101001011: io_out <= 8'b00001000;
        11'b10101001100: io_out <= 8'b00001000;
        11'b10101001101: io_out <= 8'b00001000;
        11'b10101001110: io_out <= 8'b00001000;
        11'b10101010001: io_out <= 8'b00001000;
        11'b10101010010: io_out <= 8'b00001000;
        11'b10101010011: io_out <= 8'b00001000;
        11'b10101010100: io_out <= 8'b00001000;
        11'b10101010101: io_out <= 8'b00001000;
        11'b10101010110: io_out <= 8'b00111000;
        11'b10101011000: io_out <= 8'b01001010;
        11'b10101011001: io_out <= 8'b00101111;
        11'b10101011010: io_out <= 8'b00011000;
        11'b10101011011: io_out <= 8'b10001000;
        11'b10101011100: io_out <= 8'b11010100;
        11'b10101011101: io_out <= 8'b11001010;
        11'b10101011110: io_out <= 8'b10101001;
        11'b10101011111: io_out <= 8'b10110000;
        11'b10101100000: io_out <= 8'b01001010;
        11'b10101100001: io_out <= 8'b00101111;
        11'b10101100010: io_out <= 8'b00011000;
        11'b10101100011: io_out <= 8'b00101000;
        11'b10101100100: io_out <= 8'b00110100;
        11'b10101100101: io_out <= 8'b00101010;
        11'b10101100110: io_out <= 8'b11111101;
        11'b10101100111: io_out <= 8'b00100000;
        11'b10101101011: io_out <= 8'b01111010;
        11'b10101110001: io_out <= 8'b00001000;
        11'b10101110010: io_out <= 8'b00010100;
        11'b10101110011: io_out <= 8'b00100010;
        11'b10101110100: io_out <= 8'b00001000;
        11'b10101110101: io_out <= 8'b00010100;
        11'b10101110110: io_out <= 8'b00100010;
        11'b10101111001: io_out <= 8'b00100010;
        11'b10101111010: io_out <= 8'b00010100;
        11'b10101111011: io_out <= 8'b00001000;
        11'b10101111100: io_out <= 8'b00100010;
        11'b10101111101: io_out <= 8'b00010100;
        11'b10101111110: io_out <= 8'b00001000;
        11'b10110000000: io_out <= 8'b10101010;
        11'b10110000010: io_out <= 8'b01010101;
        11'b10110000100: io_out <= 8'b10101010;
        11'b10110000110: io_out <= 8'b01010101;
        11'b10110001000: io_out <= 8'b10101010;
        11'b10110001001: io_out <= 8'b01010101;
        11'b10110001010: io_out <= 8'b10101010;
        11'b10110001011: io_out <= 8'b01010101;
        11'b10110001100: io_out <= 8'b10101010;
        11'b10110001101: io_out <= 8'b01010101;
        11'b10110001110: io_out <= 8'b10101010;
        11'b10110001111: io_out <= 8'b01010101;
        11'b10110010000: io_out <= 8'b11011101;
        11'b10110010001: io_out <= 8'b11111111;
        11'b10110010010: io_out <= 8'b10101010;
        11'b10110010011: io_out <= 8'b01110111;
        11'b10110010100: io_out <= 8'b11011101;
        11'b10110010101: io_out <= 8'b10101010;
        11'b10110010110: io_out <= 8'b11111111;
        11'b10110010111: io_out <= 8'b01110111;
        11'b10110011011: io_out <= 8'b11111111;
        11'b10110100000: io_out <= 8'b00010000;
        11'b10110100001: io_out <= 8'b00010000;
        11'b10110100010: io_out <= 8'b00010000;
        11'b10110100011: io_out <= 8'b11111111;
        11'b10110101000: io_out <= 8'b00010100;
        11'b10110101001: io_out <= 8'b00010100;
        11'b10110101010: io_out <= 8'b00010100;
        11'b10110101011: io_out <= 8'b11111111;
        11'b10110110000: io_out <= 8'b00010000;
        11'b10110110001: io_out <= 8'b00010000;
        11'b10110110010: io_out <= 8'b00010000;
        11'b10110110011: io_out <= 8'b11111111;
        11'b10110110101: io_out <= 8'b11111111;
        11'b10110111000: io_out <= 8'b00010000;
        11'b10110111001: io_out <= 8'b00010000;
        11'b10110111010: io_out <= 8'b00010000;
        11'b10110111011: io_out <= 8'b11110000;
        11'b10110111100: io_out <= 8'b00010000;
        11'b10110111101: io_out <= 8'b11110000;
        11'b10111000000: io_out <= 8'b00010100;
        11'b10111000001: io_out <= 8'b00010100;
        11'b10111000010: io_out <= 8'b00010100;
        11'b10111000011: io_out <= 8'b11111100;
        11'b10111001000: io_out <= 8'b00010100;
        11'b10111001001: io_out <= 8'b00010100;
        11'b10111001010: io_out <= 8'b00010100;
        11'b10111001011: io_out <= 8'b11110111;
        11'b10111001101: io_out <= 8'b11111111;
        11'b10111010011: io_out <= 8'b11111111;
        11'b10111010101: io_out <= 8'b11111111;
        11'b10111011000: io_out <= 8'b00010100;
        11'b10111011001: io_out <= 8'b00010100;
        11'b10111011010: io_out <= 8'b00010100;
        11'b10111011011: io_out <= 8'b11110100;
        11'b10111011100: io_out <= 8'b00000100;
        11'b10111011101: io_out <= 8'b11111100;
        11'b10111100000: io_out <= 8'b00010100;
        11'b10111100001: io_out <= 8'b00010100;
        11'b10111100010: io_out <= 8'b00010100;
        11'b10111100011: io_out <= 8'b00010111;
        11'b10111100100: io_out <= 8'b00010000;
        11'b10111100101: io_out <= 8'b00011111;
        11'b10111101000: io_out <= 8'b00010000;
        11'b10111101001: io_out <= 8'b00010000;
        11'b10111101010: io_out <= 8'b00010000;
        11'b10111101011: io_out <= 8'b00011111;
        11'b10111101100: io_out <= 8'b00010000;
        11'b10111101101: io_out <= 8'b00011111;
        11'b10111110000: io_out <= 8'b00010100;
        11'b10111110001: io_out <= 8'b00010100;
        11'b10111110010: io_out <= 8'b00010100;
        11'b10111110011: io_out <= 8'b00011111;
        11'b10111111000: io_out <= 8'b00010000;
        11'b10111111001: io_out <= 8'b00010000;
        11'b10111111010: io_out <= 8'b00010000;
        11'b10111111011: io_out <= 8'b11110000;
        11'b11000000011: io_out <= 8'b00011111;
        11'b11000000100: io_out <= 8'b00010000;
        11'b11000000101: io_out <= 8'b00010000;
        11'b11000000110: io_out <= 8'b00010000;
        11'b11000000111: io_out <= 8'b00010000;
        11'b11000001000: io_out <= 8'b00010000;
        11'b11000001001: io_out <= 8'b00010000;
        11'b11000001010: io_out <= 8'b00010000;
        11'b11000001011: io_out <= 8'b00011111;
        11'b11000001100: io_out <= 8'b00010000;
        11'b11000001101: io_out <= 8'b00010000;
        11'b11000001110: io_out <= 8'b00010000;
        11'b11000001111: io_out <= 8'b00010000;
        11'b11000010000: io_out <= 8'b00010000;
        11'b11000010001: io_out <= 8'b00010000;
        11'b11000010010: io_out <= 8'b00010000;
        11'b11000010011: io_out <= 8'b11110000;
        11'b11000010100: io_out <= 8'b00010000;
        11'b11000010101: io_out <= 8'b00010000;
        11'b11000010110: io_out <= 8'b00010000;
        11'b11000010111: io_out <= 8'b00010000;
        11'b11000011011: io_out <= 8'b11111111;
        11'b11000011100: io_out <= 8'b00010000;
        11'b11000011101: io_out <= 8'b00010000;
        11'b11000011110: io_out <= 8'b00010000;
        11'b11000011111: io_out <= 8'b00010000;
        11'b11000100000: io_out <= 8'b00010000;
        11'b11000100001: io_out <= 8'b00010000;
        11'b11000100010: io_out <= 8'b00010000;
        11'b11000100011: io_out <= 8'b00010000;
        11'b11000100100: io_out <= 8'b00010000;
        11'b11000100101: io_out <= 8'b00010000;
        11'b11000100110: io_out <= 8'b00010000;
        11'b11000100111: io_out <= 8'b00010000;
        11'b11000101000: io_out <= 8'b00010000;
        11'b11000101001: io_out <= 8'b00010000;
        11'b11000101010: io_out <= 8'b00010000;
        11'b11000101011: io_out <= 8'b11111111;
        11'b11000101100: io_out <= 8'b00010000;
        11'b11000101101: io_out <= 8'b00010000;
        11'b11000101110: io_out <= 8'b00010000;
        11'b11000101111: io_out <= 8'b00010000;
        11'b11000110011: io_out <= 8'b11111111;
        11'b11000110100: io_out <= 8'b00010100;
        11'b11000110101: io_out <= 8'b00010100;
        11'b11000110110: io_out <= 8'b00010100;
        11'b11000110111: io_out <= 8'b00010100;
        11'b11000111011: io_out <= 8'b11111111;
        11'b11000111101: io_out <= 8'b11111111;
        11'b11000111110: io_out <= 8'b00010000;
        11'b11000111111: io_out <= 8'b00010000;
        11'b11001000011: io_out <= 8'b00011111;
        11'b11001000100: io_out <= 8'b00010000;
        11'b11001000101: io_out <= 8'b00010111;
        11'b11001000110: io_out <= 8'b00010100;
        11'b11001000111: io_out <= 8'b00010100;
        11'b11001001011: io_out <= 8'b11111100;
        11'b11001001100: io_out <= 8'b00000100;
        11'b11001001101: io_out <= 8'b11110100;
        11'b11001001110: io_out <= 8'b00010100;
        11'b11001001111: io_out <= 8'b00010100;
        11'b11001010000: io_out <= 8'b00010100;
        11'b11001010001: io_out <= 8'b00010100;
        11'b11001010010: io_out <= 8'b00010100;
        11'b11001010011: io_out <= 8'b00010111;
        11'b11001010100: io_out <= 8'b00010000;
        11'b11001010101: io_out <= 8'b00010111;
        11'b11001010110: io_out <= 8'b00010100;
        11'b11001010111: io_out <= 8'b00010100;
        11'b11001011000: io_out <= 8'b00010100;
        11'b11001011001: io_out <= 8'b00010100;
        11'b11001011010: io_out <= 8'b00010100;
        11'b11001011011: io_out <= 8'b11110100;
        11'b11001011100: io_out <= 8'b00000100;
        11'b11001011101: io_out <= 8'b11110100;
        11'b11001011110: io_out <= 8'b00010100;
        11'b11001011111: io_out <= 8'b00010100;
        11'b11001100011: io_out <= 8'b11111111;
        11'b11001100101: io_out <= 8'b11110111;
        11'b11001100110: io_out <= 8'b00010100;
        11'b11001100111: io_out <= 8'b00010100;
        11'b11001101000: io_out <= 8'b00010100;
        11'b11001101001: io_out <= 8'b00010100;
        11'b11001101010: io_out <= 8'b00010100;
        11'b11001101011: io_out <= 8'b00010100;
        11'b11001101100: io_out <= 8'b00010100;
        11'b11001101101: io_out <= 8'b00010100;
        11'b11001101110: io_out <= 8'b00010100;
        11'b11001101111: io_out <= 8'b00010100;
        11'b11001110000: io_out <= 8'b00010100;
        11'b11001110001: io_out <= 8'b00010100;
        11'b11001110010: io_out <= 8'b00010100;
        11'b11001110011: io_out <= 8'b11110111;
        11'b11001110101: io_out <= 8'b11110111;
        11'b11001110110: io_out <= 8'b00010100;
        11'b11001110111: io_out <= 8'b00010100;
        11'b11001111000: io_out <= 8'b00010100;
        11'b11001111001: io_out <= 8'b00010100;
        11'b11001111010: io_out <= 8'b00010100;
        11'b11001111011: io_out <= 8'b00010111;
        11'b11001111100: io_out <= 8'b00010100;
        11'b11001111101: io_out <= 8'b00010100;
        11'b11001111110: io_out <= 8'b00010100;
        11'b11001111111: io_out <= 8'b00010100;
        11'b11010000000: io_out <= 8'b00010000;
        11'b11010000001: io_out <= 8'b00010000;
        11'b11010000010: io_out <= 8'b00010000;
        11'b11010000011: io_out <= 8'b00011111;
        11'b11010000100: io_out <= 8'b00010000;
        11'b11010000101: io_out <= 8'b00011111;
        11'b11010000110: io_out <= 8'b00010000;
        11'b11010000111: io_out <= 8'b00010000;
        11'b11010001000: io_out <= 8'b00010100;
        11'b11010001001: io_out <= 8'b00010100;
        11'b11010001010: io_out <= 8'b00010100;
        11'b11010001011: io_out <= 8'b11110100;
        11'b11010001100: io_out <= 8'b00010100;
        11'b11010001101: io_out <= 8'b00010100;
        11'b11010001110: io_out <= 8'b00010100;
        11'b11010001111: io_out <= 8'b00010100;
        11'b11010010000: io_out <= 8'b00010000;
        11'b11010010001: io_out <= 8'b00010000;
        11'b11010010010: io_out <= 8'b00010000;
        11'b11010010011: io_out <= 8'b11110000;
        11'b11010010100: io_out <= 8'b00010000;
        11'b11010010101: io_out <= 8'b11110000;
        11'b11010010110: io_out <= 8'b00010000;
        11'b11010010111: io_out <= 8'b00010000;
        11'b11010011011: io_out <= 8'b00011111;
        11'b11010011100: io_out <= 8'b00010000;
        11'b11010011101: io_out <= 8'b00011111;
        11'b11010011110: io_out <= 8'b00010000;
        11'b11010011111: io_out <= 8'b00010000;
        11'b11010100011: io_out <= 8'b00011111;
        11'b11010100100: io_out <= 8'b00010100;
        11'b11010100101: io_out <= 8'b00010100;
        11'b11010100110: io_out <= 8'b00010100;
        11'b11010100111: io_out <= 8'b00010100;
        11'b11010101011: io_out <= 8'b11111100;
        11'b11010101100: io_out <= 8'b00010100;
        11'b11010101101: io_out <= 8'b00010100;
        11'b11010101110: io_out <= 8'b00010100;
        11'b11010101111: io_out <= 8'b00010100;
        11'b11010110011: io_out <= 8'b11110000;
        11'b11010110100: io_out <= 8'b00010000;
        11'b11010110101: io_out <= 8'b11110000;
        11'b11010110110: io_out <= 8'b00010000;
        11'b11010110111: io_out <= 8'b00010000;
        11'b11010111000: io_out <= 8'b00010000;
        11'b11010111001: io_out <= 8'b00010000;
        11'b11010111010: io_out <= 8'b00010000;
        11'b11010111011: io_out <= 8'b11111111;
        11'b11010111100: io_out <= 8'b00010000;
        11'b11010111101: io_out <= 8'b11111111;
        11'b11010111110: io_out <= 8'b00010000;
        11'b11010111111: io_out <= 8'b00010000;
        11'b11011000000: io_out <= 8'b00010100;
        11'b11011000001: io_out <= 8'b00010100;
        11'b11011000010: io_out <= 8'b00010100;
        11'b11011000011: io_out <= 8'b11111111;
        11'b11011000100: io_out <= 8'b00010100;
        11'b11011000101: io_out <= 8'b00010100;
        11'b11011000110: io_out <= 8'b00010100;
        11'b11011000111: io_out <= 8'b00010100;
        11'b11011001000: io_out <= 8'b00010000;
        11'b11011001001: io_out <= 8'b00010000;
        11'b11011001010: io_out <= 8'b00010000;
        11'b11011001011: io_out <= 8'b00011111;
        11'b11011010011: io_out <= 8'b11110000;
        11'b11011010100: io_out <= 8'b00010000;
        11'b11011010101: io_out <= 8'b00010000;
        11'b11011010110: io_out <= 8'b00010000;
        11'b11011010111: io_out <= 8'b00010000;
        11'b11011011000: io_out <= 8'b11111111;
        11'b11011011001: io_out <= 8'b11111111;
        11'b11011011010: io_out <= 8'b11111111;
        11'b11011011011: io_out <= 8'b11111111;
        11'b11011011100: io_out <= 8'b11111111;
        11'b11011011101: io_out <= 8'b11111111;
        11'b11011011110: io_out <= 8'b11111111;
        11'b11011011111: io_out <= 8'b11111111;
        11'b11011100000: io_out <= 8'b11110000;
        11'b11011100001: io_out <= 8'b11110000;
        11'b11011100010: io_out <= 8'b11110000;
        11'b11011100011: io_out <= 8'b11110000;
        11'b11011100100: io_out <= 8'b11110000;
        11'b11011100101: io_out <= 8'b11110000;
        11'b11011100110: io_out <= 8'b11110000;
        11'b11011100111: io_out <= 8'b11110000;
        11'b11011101000: io_out <= 8'b11111111;
        11'b11011101001: io_out <= 8'b11111111;
        11'b11011101010: io_out <= 8'b11111111;
        11'b11011101011: io_out <= 8'b11111111;
        11'b11011110100: io_out <= 8'b11111111;
        11'b11011110101: io_out <= 8'b11111111;
        11'b11011110110: io_out <= 8'b11111111;
        11'b11011110111: io_out <= 8'b11111111;
        11'b11011111000: io_out <= 8'b00001111;
        11'b11011111001: io_out <= 8'b00001111;
        11'b11011111010: io_out <= 8'b00001111;
        11'b11011111011: io_out <= 8'b00001111;
        11'b11011111100: io_out <= 8'b00001111;
        11'b11011111101: io_out <= 8'b00001111;
        11'b11011111110: io_out <= 8'b00001111;
        11'b11011111111: io_out <= 8'b00001111;
        11'b11100000001: io_out <= 8'b00111000;
        11'b11100000010: io_out <= 8'b01000100;
        11'b11100000011: io_out <= 8'b01000100;
        11'b11100000100: io_out <= 8'b00101000;
        11'b11100000101: io_out <= 8'b00010000;
        11'b11100000110: io_out <= 8'b00101000;
        11'b11100000111: io_out <= 8'b01000100;
        11'b11100001001: io_out <= 8'b11111100;
        11'b11100001010: io_out <= 8'b00101010;
        11'b11100001011: io_out <= 8'b00101010;
        11'b11100001100: io_out <= 8'b00101010;
        11'b11100001101: io_out <= 8'b00101010;
        11'b11100001110: io_out <= 8'b00010100;
        11'b11100010001: io_out <= 8'b01111110;
        11'b11100010010: io_out <= 8'b00000010;
        11'b11100010011: io_out <= 8'b00000010;
        11'b11100010100: io_out <= 8'b00000010;
        11'b11100010101: io_out <= 8'b00000010;
        11'b11100010110: io_out <= 8'b00000110;
        11'b11100011001: io_out <= 8'b00000100;
        11'b11100011010: io_out <= 8'b00000010;
        11'b11100011011: io_out <= 8'b01111110;
        11'b11100011100: io_out <= 8'b00000010;
        11'b11100011101: io_out <= 8'b01111110;
        11'b11100011110: io_out <= 8'b00000010;
        11'b11100011111: io_out <= 8'b00000010;
        11'b11100100001: io_out <= 8'b01100011;
        11'b11100100010: io_out <= 8'b01010101;
        11'b11100100011: io_out <= 8'b01001001;
        11'b11100100100: io_out <= 8'b01001001;
        11'b11100100101: io_out <= 8'b01000001;
        11'b11100100110: io_out <= 8'b01100011;
        11'b11100101001: io_out <= 8'b00111000;
        11'b11100101010: io_out <= 8'b01000100;
        11'b11100101011: io_out <= 8'b01000100;
        11'b11100101100: io_out <= 8'b00111100;
        11'b11100101101: io_out <= 8'b00000100;
        11'b11100101110: io_out <= 8'b00000100;
        11'b11100110000: io_out <= 8'b10000000;
        11'b11100110001: io_out <= 8'b01111110;
        11'b11100110010: io_out <= 8'b00010000;
        11'b11100110011: io_out <= 8'b00010000;
        11'b11100110100: io_out <= 8'b00010000;
        11'b11100110101: io_out <= 8'b00001110;
        11'b11100110110: io_out <= 8'b00010000;
        11'b11100111001: io_out <= 8'b00000100;
        11'b11100111010: io_out <= 8'b00000010;
        11'b11100111011: io_out <= 8'b00000010;
        11'b11100111100: io_out <= 8'b01111100;
        11'b11100111101: io_out <= 8'b00000100;
        11'b11100111110: io_out <= 8'b00000010;
        11'b11100111111: io_out <= 8'b00000010;
        11'b11101000001: io_out <= 8'b10011001;
        11'b11101000010: io_out <= 8'b10100101;
        11'b11101000011: io_out <= 8'b11100111;
        11'b11101000100: io_out <= 8'b10100101;
        11'b11101000101: io_out <= 8'b10011001;
        11'b11101001001: io_out <= 8'b00011100;
        11'b11101001010: io_out <= 8'b00101010;
        11'b11101001011: io_out <= 8'b01001001;
        11'b11101001100: io_out <= 8'b01001001;
        11'b11101001101: io_out <= 8'b00101010;
        11'b11101001110: io_out <= 8'b00011100;
        11'b11101010001: io_out <= 8'b01001100;
        11'b11101010010: io_out <= 8'b01110010;
        11'b11101010011: io_out <= 8'b00000001;
        11'b11101010100: io_out <= 8'b00000001;
        11'b11101010101: io_out <= 8'b01110010;
        11'b11101010110: io_out <= 8'b01001100;
        11'b11101011001: io_out <= 8'b00110000;
        11'b11101011010: io_out <= 8'b01001010;
        11'b11101011011: io_out <= 8'b01001101;
        11'b11101011100: io_out <= 8'b01001101;
        11'b11101011101: io_out <= 8'b01001001;
        11'b11101011110: io_out <= 8'b00110000;
        11'b11101100000: io_out <= 8'b00011100;
        11'b11101100001: io_out <= 8'b00100010;
        11'b11101100010: io_out <= 8'b00100010;
        11'b11101100011: io_out <= 8'b00010100;
        11'b11101100100: io_out <= 8'b00001000;
        11'b11101100101: io_out <= 8'b00010100;
        11'b11101100110: io_out <= 8'b00100010;
        11'b11101100111: io_out <= 8'b00011100;
        11'b11101101000: io_out <= 8'b10000000;
        11'b11101101001: io_out <= 8'b01011000;
        11'b11101101010: io_out <= 8'b00100100;
        11'b11101101011: io_out <= 8'b00110100;
        11'b11101101100: io_out <= 8'b00101100;
        11'b11101101101: io_out <= 8'b00100110;
        11'b11101101110: io_out <= 8'b00011001;
        11'b11101110010: io_out <= 8'b00011100;
        11'b11101110011: io_out <= 8'b00101010;
        11'b11101110100: io_out <= 8'b01001001;
        11'b11101110101: io_out <= 8'b01001001;
        11'b11101111001: io_out <= 8'b01111110;
        11'b11101111010: io_out <= 8'b00000001;
        11'b11101111011: io_out <= 8'b00000001;
        11'b11101111100: io_out <= 8'b00000001;
        11'b11101111101: io_out <= 8'b00000001;
        11'b11101111110: io_out <= 8'b01111110;
        11'b11110000001: io_out <= 8'b00101010;
        11'b11110000010: io_out <= 8'b00101010;
        11'b11110000011: io_out <= 8'b00101010;
        11'b11110000100: io_out <= 8'b00101010;
        11'b11110000101: io_out <= 8'b00101010;
        11'b11110000110: io_out <= 8'b00101010;
        11'b11110001001: io_out <= 8'b01000100;
        11'b11110001010: io_out <= 8'b01000100;
        11'b11110001011: io_out <= 8'b01011111;
        11'b11110001100: io_out <= 8'b01000100;
        11'b11110001101: io_out <= 8'b01000100;
        11'b11110010001: io_out <= 8'b01000000;
        11'b11110010010: io_out <= 8'b01000000;
        11'b11110010011: io_out <= 8'b01010001;
        11'b11110010100: io_out <= 8'b01001010;
        11'b11110010101: io_out <= 8'b01000100;
        11'b11110010110: io_out <= 8'b01000000;
        11'b11110011001: io_out <= 8'b01000000;
        11'b11110011010: io_out <= 8'b01000100;
        11'b11110011011: io_out <= 8'b01001010;
        11'b11110011100: io_out <= 8'b01010001;
        11'b11110011101: io_out <= 8'b01000000;
        11'b11110011110: io_out <= 8'b01000000;
        11'b11110100011: io_out <= 8'b11111110;
        11'b11110100100: io_out <= 8'b00000001;
        11'b11110100101: io_out <= 8'b00000001;
        11'b11110100110: io_out <= 8'b00000110;
        11'b11110101000: io_out <= 8'b01100000;
        11'b11110101001: io_out <= 8'b10000000;
        11'b11110101010: io_out <= 8'b10000000;
        11'b11110101011: io_out <= 8'b01111111;
        11'b11110110001: io_out <= 8'b00001000;
        11'b11110110010: io_out <= 8'b00001000;
        11'b11110110011: io_out <= 8'b01101011;
        11'b11110110100: io_out <= 8'b01101011;
        11'b11110110101: io_out <= 8'b00001000;
        11'b11110110110: io_out <= 8'b00001000;
        11'b11110111001: io_out <= 8'b00100100;
        11'b11110111010: io_out <= 8'b00010010;
        11'b11110111011: io_out <= 8'b00010010;
        11'b11110111100: io_out <= 8'b00100100;
        11'b11110111101: io_out <= 8'b00100100;
        11'b11110111110: io_out <= 8'b00010010;
        11'b11111000001: io_out <= 8'b00000110;
        11'b11111000010: io_out <= 8'b00001001;
        11'b11111000011: io_out <= 8'b00001001;
        11'b11111000100: io_out <= 8'b00000110;
        11'b11111001011: io_out <= 8'b00011000;
        11'b11111001100: io_out <= 8'b00011000;
        11'b11111010011: io_out <= 8'b00010000;
        11'b11111010100: io_out <= 8'b00010000;
        11'b11111011000: io_out <= 8'b00100000;
        11'b11111011001: io_out <= 8'b00100000;
        11'b11111011010: io_out <= 8'b01000000;
        11'b11111011011: io_out <= 8'b10000000;
        11'b11111011100: io_out <= 8'b11111111;
        11'b11111011101: io_out <= 8'b00000001;
        11'b11111011110: io_out <= 8'b00000001;
        11'b11111011111: io_out <= 8'b00000001;
        11'b11111100001: io_out <= 8'b00011111;
        11'b11111100010: io_out <= 8'b00000001;
        11'b11111100011: io_out <= 8'b00000001;
        11'b11111100100: io_out <= 8'b00000001;
        11'b11111100101: io_out <= 8'b00011110;
        11'b11111101001: io_out <= 8'b00010010;
        11'b11111101010: io_out <= 8'b00011001;
        11'b11111101011: io_out <= 8'b00010101;
        11'b11111101100: io_out <= 8'b00010010;
        11'b11111110010: io_out <= 8'b00111100;
        11'b11111110011: io_out <= 8'b00111100;
        11'b11111110100: io_out <= 8'b00111100;
        11'b11111110101: io_out <= 8'b00111100;
        default: io_out <= 8'b00000000;
    endcase;
end

endmodule
